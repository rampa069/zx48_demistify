library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"0487da01",
     1 => x"580e87dd",
     2 => x"0e5a595e",
     3 => x"00002927",
     4 => x"4a260f00",
     5 => x"48264926",
     6 => x"082680ff",
     7 => x"002d274f",
     8 => x"274f0000",
     9 => x"0000002a",
    10 => x"fd004f4f",
    11 => x"d0c1c387",
    12 => x"48c0c84e",
    13 => x"d5c128c2",
    14 => x"ead6e5ea",
    15 => x"c1467149",
    16 => x"87f90188",
    17 => x"49d0c1c3",
    18 => x"48ece9c2",
    19 => x"0389d089",
    20 => x"404040c0",
    21 => x"d087f640",
    22 => x"50c00581",
    23 => x"f90589c1",
    24 => x"ece9c287",
    25 => x"e8e9c24d",
    26 => x"02ad744c",
    27 => x"0f2487c4",
    28 => x"efc187f7",
    29 => x"e9c287e6",
    30 => x"e9c24dec",
    31 => x"ad744cec",
    32 => x"c487c602",
    33 => x"f50f6c8c",
    34 => x"87fd0087",
    35 => x"7186fc1e",
    36 => x"49c0ff4a",
    37 => x"c0c44869",
    38 => x"487e7098",
    39 => x"87f40298",
    40 => x"fc487972",
    41 => x"0e4f268e",
    42 => x"0e5c5b5e",
    43 => x"4cc04b71",
    44 => x"029a4a13",
    45 => x"497287cd",
    46 => x"c187d1ff",
    47 => x"9a4a1384",
    48 => x"7487f305",
    49 => x"264c2648",
    50 => x"1e4f264b",
    51 => x"1e731e72",
    52 => x"02114812",
    53 => x"c34b87ca",
    54 => x"739b98df",
    55 => x"87f00288",
    56 => x"4a264b26",
    57 => x"731e4f26",
    58 => x"c11e721e",
    59 => x"87ca048b",
    60 => x"02114812",
    61 => x"028887c4",
    62 => x"4a2687f1",
    63 => x"4f264b26",
    64 => x"731e741e",
    65 => x"c11e721e",
    66 => x"87d0048b",
    67 => x"02114812",
    68 => x"c34c87ca",
    69 => x"749c98df",
    70 => x"87eb0288",
    71 => x"4b264a26",
    72 => x"4f264c26",
    73 => x"8148731e",
    74 => x"c502a973",
    75 => x"05531287",
    76 => x"4f2687f6",
    77 => x"721e731e",
    78 => x"e7c0029a",
    79 => x"c148c087",
    80 => x"06a9724b",
    81 => x"827287d1",
    82 => x"7387c906",
    83 => x"01a97283",
    84 => x"87c387f4",
    85 => x"723ab2c1",
    86 => x"738903a9",
    87 => x"2ac10780",
    88 => x"87f3052b",
    89 => x"4f264b26",
    90 => x"c41e751e",
    91 => x"a1b7714d",
    92 => x"c1b9ff04",
    93 => x"07bdc381",
    94 => x"04a2b772",
    95 => x"82c1baff",
    96 => x"fe07bdc1",
    97 => x"2dc187ee",
    98 => x"c1b8ff04",
    99 => x"042d0780",
   100 => x"81c1b9ff",
   101 => x"264d2607",
   102 => x"1e731e4f",
   103 => x"66c84a71",
   104 => x"8bc1494b",
   105 => x"cf029971",
   106 => x"ff481287",
   107 => x"737808d4",
   108 => x"718bc149",
   109 => x"87f10599",
   110 => x"4f264b26",
   111 => x"5c5b5e0e",
   112 => x"ff4a710e",
   113 => x"66cc4cd4",
   114 => x"8bc1494b",
   115 => x"ce029971",
   116 => x"7cffc387",
   117 => x"4973526c",
   118 => x"99718bc1",
   119 => x"2687f205",
   120 => x"264b264c",
   121 => x"1e731e4f",
   122 => x"c34bd4ff",
   123 => x"4a6b7bff",
   124 => x"6b7bffc3",
   125 => x"7232c849",
   126 => x"7bffc3b1",
   127 => x"31c84a6b",
   128 => x"ffc3b271",
   129 => x"c8496b7b",
   130 => x"71b17232",
   131 => x"264b2648",
   132 => x"5b5e0e4f",
   133 => x"710e5d5c",
   134 => x"4cd4ff4d",
   135 => x"ffc34875",
   136 => x"c27c7098",
   137 => x"05bfece9",
   138 => x"66d087c8",
   139 => x"d430c948",
   140 => x"66d058a6",
   141 => x"7129d849",
   142 => x"98ffc348",
   143 => x"66d07c70",
   144 => x"7129d049",
   145 => x"98ffc348",
   146 => x"66d07c70",
   147 => x"7129c849",
   148 => x"98ffc348",
   149 => x"66d07c70",
   150 => x"98ffc348",
   151 => x"49757c70",
   152 => x"487129d0",
   153 => x"7098ffc3",
   154 => x"c94b6c7c",
   155 => x"c34afff0",
   156 => x"cf05abff",
   157 => x"7c714987",
   158 => x"8ac14b6c",
   159 => x"7187c502",
   160 => x"87f202ab",
   161 => x"4d264873",
   162 => x"4b264c26",
   163 => x"c01e4f26",
   164 => x"48d4ff49",
   165 => x"c178ffc3",
   166 => x"b7c8c381",
   167 => x"87f104a9",
   168 => x"5e0e4f26",
   169 => x"0e5d5c5b",
   170 => x"c1f0ffc0",
   171 => x"c0c14df7",
   172 => x"c0c0c0c0",
   173 => x"87d6ff4b",
   174 => x"4cdff8c4",
   175 => x"49751ec0",
   176 => x"c487cefd",
   177 => x"05a8c186",
   178 => x"ff87e5c0",
   179 => x"ffc348d4",
   180 => x"c01e7378",
   181 => x"e9c1f0e1",
   182 => x"87f5fc49",
   183 => x"987086c4",
   184 => x"ff87ca05",
   185 => x"ffc348d4",
   186 => x"cb48c178",
   187 => x"87defe87",
   188 => x"ff058cc1",
   189 => x"48c087c6",
   190 => x"4c264d26",
   191 => x"4f264b26",
   192 => x"5c5b5e0e",
   193 => x"f0ffc00e",
   194 => x"ff4cc1c1",
   195 => x"ffc348d4",
   196 => x"49c4cd78",
   197 => x"d387d0f6",
   198 => x"741ec04b",
   199 => x"87f1fb49",
   200 => x"987086c4",
   201 => x"ff87ca05",
   202 => x"ffc348d4",
   203 => x"cb48c178",
   204 => x"87dafd87",
   205 => x"ff058bc1",
   206 => x"48c087df",
   207 => x"4b264c26",
   208 => x"00004f26",
   209 => x"00444d43",
   210 => x"5c5b5e0e",
   211 => x"ffc30e5d",
   212 => x"4bd4ff4d",
   213 => x"c687f7fc",
   214 => x"e1c01eea",
   215 => x"49c8c1f0",
   216 => x"c487eefa",
   217 => x"02a8c186",
   218 => x"d3fe87c8",
   219 => x"c148c087",
   220 => x"f0f987e8",
   221 => x"cf497087",
   222 => x"c699ffff",
   223 => x"c802a9ea",
   224 => x"87fcfd87",
   225 => x"d1c148c0",
   226 => x"c07b7587",
   227 => x"d1fc4cf1",
   228 => x"02987087",
   229 => x"c087ecc0",
   230 => x"f0ffc01e",
   231 => x"f949fac1",
   232 => x"86c487ef",
   233 => x"da059870",
   234 => x"6b7b7587",
   235 => x"757b7549",
   236 => x"757b757b",
   237 => x"99c0c17b",
   238 => x"c187c402",
   239 => x"c087db48",
   240 => x"c287d748",
   241 => x"87ca05ac",
   242 => x"f349e4cf",
   243 => x"48c087d9",
   244 => x"8cc187c8",
   245 => x"87f6fe05",
   246 => x"4d2648c0",
   247 => x"4b264c26",
   248 => x"00004f26",
   249 => x"43484453",
   250 => x"69616620",
   251 => x"000a216c",
   252 => x"5c5b5e0e",
   253 => x"d0ff0e5d",
   254 => x"d0e5c04d",
   255 => x"c24cc0c1",
   256 => x"c148ece9",
   257 => x"49fcd178",
   258 => x"c787dcf2",
   259 => x"f97dc24b",
   260 => x"7dc387fc",
   261 => x"49741ec0",
   262 => x"c487f6f7",
   263 => x"05a8c186",
   264 => x"c24b87c1",
   265 => x"87cb05ab",
   266 => x"f149f4d1",
   267 => x"48c087f9",
   268 => x"c187f6c0",
   269 => x"d4ff058b",
   270 => x"87ccfc87",
   271 => x"58f0e9c2",
   272 => x"cd059870",
   273 => x"c01ec187",
   274 => x"d0c1f0ff",
   275 => x"87c1f749",
   276 => x"d4ff86c4",
   277 => x"78ffc348",
   278 => x"c287ccc5",
   279 => x"c258f4e9",
   280 => x"48d4ff7d",
   281 => x"c178ffc3",
   282 => x"264d2648",
   283 => x"264b264c",
   284 => x"0000004f",
   285 => x"52524549",
   286 => x"00000000",
   287 => x"00495053",
   288 => x"5c5b5e0e",
   289 => x"4d710e5d",
   290 => x"ff4cffc3",
   291 => x"7b744bd4",
   292 => x"c448d0ff",
   293 => x"7b7478c3",
   294 => x"ffc01e75",
   295 => x"49d8c1f0",
   296 => x"c487eef5",
   297 => x"02987086",
   298 => x"ecd387cb",
   299 => x"87f7ef49",
   300 => x"eec048c1",
   301 => x"c37b7487",
   302 => x"c0c87bfe",
   303 => x"4966d41e",
   304 => x"c487d6f3",
   305 => x"747b7486",
   306 => x"d87b747b",
   307 => x"744ae0da",
   308 => x"c5056b7b",
   309 => x"058ac187",
   310 => x"7b7487f5",
   311 => x"c248d0ff",
   312 => x"2648c078",
   313 => x"264c264d",
   314 => x"004f264b",
   315 => x"74697257",
   316 => x"61662065",
   317 => x"64656c69",
   318 => x"5e0e000a",
   319 => x"0e5d5c5b",
   320 => x"4b7186fc",
   321 => x"c04cd4ff",
   322 => x"cdeec57e",
   323 => x"ffc34adf",
   324 => x"c3486c7c",
   325 => x"c005a8fe",
   326 => x"4d7487f8",
   327 => x"cc029b73",
   328 => x"1e66d487",
   329 => x"d3f24973",
   330 => x"d486c487",
   331 => x"48d0ff87",
   332 => x"d478d1c4",
   333 => x"ffc34a66",
   334 => x"058ac17d",
   335 => x"a6d887f8",
   336 => x"7cffc35a",
   337 => x"059b737c",
   338 => x"d0ff87c5",
   339 => x"c178d048",
   340 => x"8ac17e4a",
   341 => x"87f6fe05",
   342 => x"8efc486e",
   343 => x"4c264d26",
   344 => x"4f264b26",
   345 => x"711e731e",
   346 => x"ff4bc04a",
   347 => x"ffc348d4",
   348 => x"48d0ff78",
   349 => x"ff78c3c4",
   350 => x"ffc348d4",
   351 => x"c01e7278",
   352 => x"d1c1f0ff",
   353 => x"87c9f249",
   354 => x"987086c4",
   355 => x"c887d205",
   356 => x"66cc1ec0",
   357 => x"87e2fd49",
   358 => x"4b7086c4",
   359 => x"c248d0ff",
   360 => x"26487378",
   361 => x"0e4f264b",
   362 => x"5d5c5b5e",
   363 => x"c01ec00e",
   364 => x"c9c1f0ff",
   365 => x"87d9f149",
   366 => x"e9c21ed2",
   367 => x"f9fc49f4",
   368 => x"c086c887",
   369 => x"d284c14c",
   370 => x"f804acb7",
   371 => x"f4e9c287",
   372 => x"c349bf97",
   373 => x"c0c199c0",
   374 => x"e7c005a9",
   375 => x"fbe9c287",
   376 => x"d049bf97",
   377 => x"fce9c231",
   378 => x"c84abf97",
   379 => x"c2b17232",
   380 => x"bf97fde9",
   381 => x"4c71b14a",
   382 => x"ffffffcf",
   383 => x"ca84c19c",
   384 => x"87e7c134",
   385 => x"97fde9c2",
   386 => x"31c149bf",
   387 => x"e9c299c6",
   388 => x"4abf97fe",
   389 => x"722ab7c7",
   390 => x"f9e9c2b1",
   391 => x"4d4abf97",
   392 => x"e9c29dcf",
   393 => x"4abf97fa",
   394 => x"32ca9ac3",
   395 => x"97fbe9c2",
   396 => x"33c24bbf",
   397 => x"e9c2b273",
   398 => x"4bbf97fc",
   399 => x"c69bc0c3",
   400 => x"b2732bb7",
   401 => x"48c181c2",
   402 => x"49703071",
   403 => x"307548c1",
   404 => x"4c724d70",
   405 => x"947184c1",
   406 => x"adb7c0c8",
   407 => x"c187cc06",
   408 => x"c82db734",
   409 => x"01adb7c0",
   410 => x"7487f4ff",
   411 => x"264d2648",
   412 => x"264b264c",
   413 => x"5b5e0e4f",
   414 => x"f80e5d5c",
   415 => x"dcf2c286",
   416 => x"c278c048",
   417 => x"c01ed4ea",
   418 => x"87d8fb49",
   419 => x"987086c4",
   420 => x"c087c505",
   421 => x"87c0c948",
   422 => x"7ec14dc0",
   423 => x"bff8fec0",
   424 => x"caebc249",
   425 => x"4bc8714a",
   426 => x"7087fbe8",
   427 => x"87c20598",
   428 => x"fec07ec0",
   429 => x"c249bff4",
   430 => x"714ae6eb",
   431 => x"e5e84bc8",
   432 => x"05987087",
   433 => x"7ec087c2",
   434 => x"fdc0026e",
   435 => x"daf1c287",
   436 => x"f2c24dbf",
   437 => x"7ebf9fd2",
   438 => x"ead6c548",
   439 => x"87c705a8",
   440 => x"bfdaf1c2",
   441 => x"6e87ce4d",
   442 => x"d5e9ca48",
   443 => x"87c502a8",
   444 => x"e3c748c0",
   445 => x"d4eac287",
   446 => x"f949751e",
   447 => x"86c487e6",
   448 => x"c5059870",
   449 => x"c748c087",
   450 => x"fec087ce",
   451 => x"c249bff4",
   452 => x"714ae6eb",
   453 => x"cde74bc8",
   454 => x"05987087",
   455 => x"f2c287c8",
   456 => x"78c148dc",
   457 => x"fec087da",
   458 => x"c249bff8",
   459 => x"714acaeb",
   460 => x"f1e64bc8",
   461 => x"02987087",
   462 => x"c087c5c0",
   463 => x"87d8c648",
   464 => x"97d2f2c2",
   465 => x"d5c149bf",
   466 => x"cdc005a9",
   467 => x"d3f2c287",
   468 => x"c249bf97",
   469 => x"c002a9ea",
   470 => x"48c087c5",
   471 => x"c287f9c5",
   472 => x"bf97d4ea",
   473 => x"e9c3487e",
   474 => x"cec002a8",
   475 => x"c3486e87",
   476 => x"c002a8eb",
   477 => x"48c087c5",
   478 => x"c287ddc5",
   479 => x"bf97dfea",
   480 => x"c0059949",
   481 => x"eac287cc",
   482 => x"49bf97e0",
   483 => x"c002a9c2",
   484 => x"48c087c5",
   485 => x"c287c1c5",
   486 => x"bf97e1ea",
   487 => x"d8f2c248",
   488 => x"484c7058",
   489 => x"f2c288c1",
   490 => x"eac258dc",
   491 => x"49bf97e2",
   492 => x"eac28175",
   493 => x"4abf97e3",
   494 => x"a17232c8",
   495 => x"ecf6c27e",
   496 => x"c2786e48",
   497 => x"bf97e4ea",
   498 => x"58a6c848",
   499 => x"bfdcf2c2",
   500 => x"87cfc202",
   501 => x"bff4fec0",
   502 => x"e6ebc249",
   503 => x"4bc8714a",
   504 => x"7087c3e4",
   505 => x"c5c00298",
   506 => x"c348c087",
   507 => x"f2c287ea",
   508 => x"c24cbfd4",
   509 => x"c25cc0f7",
   510 => x"bf97f9ea",
   511 => x"c231c849",
   512 => x"bf97f8ea",
   513 => x"c249a14a",
   514 => x"bf97faea",
   515 => x"7232d04a",
   516 => x"eac249a1",
   517 => x"4abf97fb",
   518 => x"a17232d8",
   519 => x"9166c449",
   520 => x"bfecf6c2",
   521 => x"f4f6c281",
   522 => x"c1ebc259",
   523 => x"c84abf97",
   524 => x"c0ebc232",
   525 => x"a24bbf97",
   526 => x"c2ebc24a",
   527 => x"d04bbf97",
   528 => x"4aa27333",
   529 => x"97c3ebc2",
   530 => x"9bcf4bbf",
   531 => x"a27333d8",
   532 => x"f8f6c24a",
   533 => x"748ac25a",
   534 => x"f8f6c292",
   535 => x"78a17248",
   536 => x"c287c1c1",
   537 => x"bf97e6ea",
   538 => x"c231c849",
   539 => x"bf97e5ea",
   540 => x"c549a14a",
   541 => x"81ffc731",
   542 => x"f7c229c9",
   543 => x"eac259c0",
   544 => x"4abf97eb",
   545 => x"eac232c8",
   546 => x"4bbf97ea",
   547 => x"66c44aa2",
   548 => x"c2826e92",
   549 => x"c25afcf6",
   550 => x"c048f4f6",
   551 => x"f0f6c278",
   552 => x"78a17248",
   553 => x"48c0f7c2",
   554 => x"bff4f6c2",
   555 => x"c4f7c278",
   556 => x"f8f6c248",
   557 => x"f2c278bf",
   558 => x"c002bfdc",
   559 => x"487487c9",
   560 => x"7e7030c4",
   561 => x"c287c9c0",
   562 => x"48bffcf6",
   563 => x"7e7030c4",
   564 => x"48e0f2c2",
   565 => x"48c1786e",
   566 => x"4d268ef8",
   567 => x"4b264c26",
   568 => x"5e0e4f26",
   569 => x"0e5d5c5b",
   570 => x"f2c24a71",
   571 => x"cb02bfdc",
   572 => x"c74b7287",
   573 => x"c14d722b",
   574 => x"87c99dff",
   575 => x"2bc84b72",
   576 => x"ffc34d72",
   577 => x"ecf6c29d",
   578 => x"fec083bf",
   579 => x"02abbff0",
   580 => x"fec087d9",
   581 => x"eac25bf4",
   582 => x"49731ed4",
   583 => x"c487c5f1",
   584 => x"05987086",
   585 => x"48c087c5",
   586 => x"c287e6c0",
   587 => x"02bfdcf2",
   588 => x"497587d2",
   589 => x"eac291c4",
   590 => x"4c6981d4",
   591 => x"ffffffcf",
   592 => x"87cb9cff",
   593 => x"91c24975",
   594 => x"81d4eac2",
   595 => x"744c699f",
   596 => x"264d2648",
   597 => x"264b264c",
   598 => x"5b5e0e4f",
   599 => x"f00e5d5c",
   600 => x"59a6cc86",
   601 => x"c50566c8",
   602 => x"c448c087",
   603 => x"66c887c4",
   604 => x"7080c848",
   605 => x"78c0487e",
   606 => x"0266e0c0",
   607 => x"e0c087c8",
   608 => x"05bf9766",
   609 => x"48c087c5",
   610 => x"c087e7c3",
   611 => x"4949c11e",
   612 => x"c487e5d0",
   613 => x"9c4c7086",
   614 => x"87fec002",
   615 => x"4ae4f2c2",
   616 => x"4966e0c0",
   617 => x"87e3dcff",
   618 => x"c0029870",
   619 => x"4a7487ec",
   620 => x"4966e0c0",
   621 => x"ddff4bcb",
   622 => x"987087c6",
   623 => x"c087db02",
   624 => x"029c741e",
   625 => x"4dc087c4",
   626 => x"4dc187c2",
   627 => x"e7cf4975",
   628 => x"7086c487",
   629 => x"ff059c4c",
   630 => x"9c7487c2",
   631 => x"87d0c202",
   632 => x"6e49a4dc",
   633 => x"da786948",
   634 => x"66c849a4",
   635 => x"c880c448",
   636 => x"699f58a6",
   637 => x"0866c448",
   638 => x"dcf2c278",
   639 => x"87d202bf",
   640 => x"9f49a4d4",
   641 => x"ffc04969",
   642 => x"487199ff",
   643 => x"58a630d0",
   644 => x"a6cc87c5",
   645 => x"cc78c048",
   646 => x"66c44866",
   647 => x"66c480bf",
   648 => x"66c87808",
   649 => x"c878c048",
   650 => x"81cc4966",
   651 => x"79bf66c4",
   652 => x"d04966c8",
   653 => x"4d79c081",
   654 => x"c84c66c4",
   655 => x"82d44a66",
   656 => x"91c84975",
   657 => x"c049a172",
   658 => x"c1796c41",
   659 => x"adb7c685",
   660 => x"87e7ff04",
   661 => x"c94abf6e",
   662 => x"c049722a",
   663 => x"dbff4af0",
   664 => x"4a7087d2",
   665 => x"c14966c8",
   666 => x"797281c4",
   667 => x"87c248c1",
   668 => x"8ef048c0",
   669 => x"4c264d26",
   670 => x"4f264b26",
   671 => x"5c5b5e0e",
   672 => x"4c710e5d",
   673 => x"744d66d0",
   674 => x"c2c1029c",
   675 => x"49a4c887",
   676 => x"fac00269",
   677 => x"85496c87",
   678 => x"f2c2b975",
   679 => x"ff4abfd8",
   680 => x"719972ba",
   681 => x"e4c00299",
   682 => x"4ba4c487",
   683 => x"f1f8496b",
   684 => x"c27b7087",
   685 => x"49bfd4f2",
   686 => x"7c71816c",
   687 => x"f2c2b975",
   688 => x"ff4abfd8",
   689 => x"719972ba",
   690 => x"dcff0599",
   691 => x"267c7587",
   692 => x"264c264d",
   693 => x"1e4f264b",
   694 => x"4b711e73",
   695 => x"87c7029b",
   696 => x"6949a3c8",
   697 => x"c087c505",
   698 => x"87f6c048",
   699 => x"bff0f6c2",
   700 => x"4aa3c449",
   701 => x"8ac24a6a",
   702 => x"bfd4f2c2",
   703 => x"49a17292",
   704 => x"bfd8f2c2",
   705 => x"729a6b4a",
   706 => x"fec049a1",
   707 => x"66c859f4",
   708 => x"cfe9711e",
   709 => x"7086c487",
   710 => x"87c40598",
   711 => x"87c248c0",
   712 => x"4b2648c1",
   713 => x"731e4f26",
   714 => x"9b4b711e",
   715 => x"c887c702",
   716 => x"056949a3",
   717 => x"48c087c5",
   718 => x"c287f6c0",
   719 => x"49bff0f6",
   720 => x"6a4aa3c4",
   721 => x"c28ac24a",
   722 => x"92bfd4f2",
   723 => x"c249a172",
   724 => x"4abfd8f2",
   725 => x"a1729a6b",
   726 => x"f4fec049",
   727 => x"1e66c859",
   728 => x"87dce471",
   729 => x"987086c4",
   730 => x"c087c405",
   731 => x"c187c248",
   732 => x"264b2648",
   733 => x"5b5e0e4f",
   734 => x"f80e5d5c",
   735 => x"c47e7186",
   736 => x"78ff48a6",
   737 => x"ffffffc1",
   738 => x"c04dffff",
   739 => x"d44a6e4b",
   740 => x"c8497382",
   741 => x"49a17291",
   742 => x"694c66d8",
   743 => x"acb7c08c",
   744 => x"7587cb04",
   745 => x"c503acb7",
   746 => x"5ba6c887",
   747 => x"83c14d74",
   748 => x"04abb7c6",
   749 => x"c487d6ff",
   750 => x"8ef84866",
   751 => x"4c264d26",
   752 => x"4f264b26",
   753 => x"5c5b5e0e",
   754 => x"86f00e5d",
   755 => x"a6c47e71",
   756 => x"ffffc148",
   757 => x"78ffffff",
   758 => x"78ff80c4",
   759 => x"4cc04dc0",
   760 => x"83d44b6e",
   761 => x"92c84a74",
   762 => x"754aa273",
   763 => x"7391c849",
   764 => x"486a49a1",
   765 => x"a6d08869",
   766 => x"02ad7458",
   767 => x"66c487cf",
   768 => x"87c903a8",
   769 => x"c45ca6cc",
   770 => x"66cc48a6",
   771 => x"c684c178",
   772 => x"ff04acb7",
   773 => x"85c187ca",
   774 => x"04adb7c6",
   775 => x"c887fffe",
   776 => x"8ef04866",
   777 => x"4c264d26",
   778 => x"4f264b26",
   779 => x"5c5b5e0e",
   780 => x"86ec0e5d",
   781 => x"e4c04b71",
   782 => x"28c94866",
   783 => x"c258a6c8",
   784 => x"4abfd8f2",
   785 => x"4872baff",
   786 => x"cc9866c4",
   787 => x"9b7358a6",
   788 => x"87c1c302",
   789 => x"6949a3c8",
   790 => x"87f9c202",
   791 => x"986b4872",
   792 => x"c458a6d4",
   793 => x"7e6c4ca3",
   794 => x"d04866c8",
   795 => x"c605a866",
   796 => x"7b66c487",
   797 => x"c887ccc2",
   798 => x"49731e66",
   799 => x"c487f6fb",
   800 => x"c04d7086",
   801 => x"d004adb7",
   802 => x"4aa3d487",
   803 => x"91c84975",
   804 => x"2149a172",
   805 => x"c77c697b",
   806 => x"cc7bc087",
   807 => x"7c6949a3",
   808 => x"6b4866c4",
   809 => x"58a6c888",
   810 => x"731e66d0",
   811 => x"87c5fb49",
   812 => x"4d7086c4",
   813 => x"49a3c4c1",
   814 => x"6948a6c8",
   815 => x"4866d078",
   816 => x"06a866c8",
   817 => x"c087f2c0",
   818 => x"c004adb7",
   819 => x"a6cc87eb",
   820 => x"78a3d448",
   821 => x"91c84975",
   822 => x"d08166cc",
   823 => x"88694866",
   824 => x"66c84970",
   825 => x"87d106a9",
   826 => x"d7fb4973",
   827 => x"c8497087",
   828 => x"8166cc91",
   829 => x"6e4166d0",
   830 => x"1e66c479",
   831 => x"fbf54973",
   832 => x"c286c487",
   833 => x"731ed4ea",
   834 => x"87cbf749",
   835 => x"a3d086c4",
   836 => x"66e4c049",
   837 => x"268eec79",
   838 => x"264c264d",
   839 => x"1e4f264b",
   840 => x"4b711e73",
   841 => x"e4c0029b",
   842 => x"c4f7c287",
   843 => x"c24a735b",
   844 => x"d4f2c28a",
   845 => x"c29249bf",
   846 => x"48bff0f6",
   847 => x"f7c28072",
   848 => x"487158c8",
   849 => x"f2c230c4",
   850 => x"edc058e4",
   851 => x"c0f7c287",
   852 => x"f4f6c248",
   853 => x"f7c278bf",
   854 => x"f6c248c4",
   855 => x"c278bff8",
   856 => x"02bfdcf2",
   857 => x"f2c287c9",
   858 => x"c449bfd4",
   859 => x"c287c731",
   860 => x"49bffcf6",
   861 => x"f2c231c4",
   862 => x"4b2659e4",
   863 => x"5e0e4f26",
   864 => x"710e5c5b",
   865 => x"724bc04a",
   866 => x"e0c0029a",
   867 => x"49a2da87",
   868 => x"c24b699f",
   869 => x"02bfdcf2",
   870 => x"a2d487cf",
   871 => x"49699f49",
   872 => x"ffffc04c",
   873 => x"c234d09c",
   874 => x"744cc087",
   875 => x"fd4973b3",
   876 => x"4c2687ed",
   877 => x"4f264b26",
   878 => x"5c5b5e0e",
   879 => x"86f00e5d",
   880 => x"cf59a6c8",
   881 => x"f8ffffff",
   882 => x"c47ec04c",
   883 => x"87d80266",
   884 => x"48d0eac2",
   885 => x"eac278c0",
   886 => x"f7c248c8",
   887 => x"c278bfc4",
   888 => x"c248ccea",
   889 => x"78bfc0f7",
   890 => x"48f1f2c2",
   891 => x"f2c250c0",
   892 => x"c249bfe0",
   893 => x"4abfd0ea",
   894 => x"c403aa71",
   895 => x"497287cc",
   896 => x"c00599cf",
   897 => x"fec087ea",
   898 => x"eac248f0",
   899 => x"c278bfc8",
   900 => x"c21ed4ea",
   901 => x"49bfc8ea",
   902 => x"48c8eac2",
   903 => x"7178a1c1",
   904 => x"87c0ddff",
   905 => x"fec086c4",
   906 => x"eac248ec",
   907 => x"87cc78d4",
   908 => x"bfecfec0",
   909 => x"80e0c048",
   910 => x"58f0fec0",
   911 => x"bfd0eac2",
   912 => x"c280c148",
   913 => x"2758d4ea",
   914 => x"00000fac",
   915 => x"4dbf97bf",
   916 => x"e5c2029d",
   917 => x"ade5c387",
   918 => x"87dec202",
   919 => x"bfecfec0",
   920 => x"49a3cb4b",
   921 => x"accf4c11",
   922 => x"87d2c105",
   923 => x"99df4975",
   924 => x"91cd89c1",
   925 => x"81e4f2c2",
   926 => x"124aa3c1",
   927 => x"4aa3c351",
   928 => x"a3c55112",
   929 => x"c751124a",
   930 => x"51124aa3",
   931 => x"124aa3c9",
   932 => x"4aa3ce51",
   933 => x"a3d05112",
   934 => x"d251124a",
   935 => x"51124aa3",
   936 => x"124aa3d4",
   937 => x"4aa3d651",
   938 => x"a3d85112",
   939 => x"dc51124a",
   940 => x"51124aa3",
   941 => x"124aa3de",
   942 => x"c07ec151",
   943 => x"497487fc",
   944 => x"c00599c8",
   945 => x"497487ed",
   946 => x"d30599d0",
   947 => x"66e0c087",
   948 => x"87ccc002",
   949 => x"e0c04973",
   950 => x"98700f66",
   951 => x"87d3c002",
   952 => x"c6c0056e",
   953 => x"e4f2c287",
   954 => x"c050c048",
   955 => x"48bfecfe",
   956 => x"c287e9c2",
   957 => x"c048f1f2",
   958 => x"f2c27e50",
   959 => x"c249bfe0",
   960 => x"4abfd0ea",
   961 => x"fb04aa71",
   962 => x"ffcf87f4",
   963 => x"4cf8ffff",
   964 => x"bfc4f7c2",
   965 => x"87c8c005",
   966 => x"bfdcf2c2",
   967 => x"87fac102",
   968 => x"bfcceac2",
   969 => x"87fae649",
   970 => x"58d0eac2",
   971 => x"c248a6c4",
   972 => x"78bfccea",
   973 => x"bfdcf2c2",
   974 => x"87dbc002",
   975 => x"744966c4",
   976 => x"02a97499",
   977 => x"c887c8c0",
   978 => x"78c048a6",
   979 => x"c887e7c0",
   980 => x"78c148a6",
   981 => x"c487dfc0",
   982 => x"ffcf4966",
   983 => x"02a999f8",
   984 => x"cc87c8c0",
   985 => x"78c048a6",
   986 => x"cc87c5c0",
   987 => x"78c148a6",
   988 => x"cc48a6c8",
   989 => x"66c87866",
   990 => x"87dec005",
   991 => x"c24966c4",
   992 => x"d4f2c289",
   993 => x"f6c291bf",
   994 => x"7148bff0",
   995 => x"cceac280",
   996 => x"d0eac258",
   997 => x"f978c048",
   998 => x"48c087d4",
   999 => x"ffffffcf",
  1000 => x"8ef04cf8",
  1001 => x"4c264d26",
  1002 => x"4f264b26",
  1003 => x"00000000",
  1004 => x"ffffffff",
  1005 => x"00000fbc",
  1006 => x"00000fc8",
  1007 => x"33544146",
  1008 => x"20202032",
  1009 => x"00000000",
  1010 => x"31544146",
  1011 => x"20202036",
  1012 => x"d4ff1e00",
  1013 => x"78ffc348",
  1014 => x"4f264868",
  1015 => x"48d4ff1e",
  1016 => x"ff78ffc3",
  1017 => x"e1c048d0",
  1018 => x"48d4ff78",
  1019 => x"4f2678d4",
  1020 => x"48d0ff1e",
  1021 => x"2678e0c0",
  1022 => x"d4ff1e4f",
  1023 => x"99497087",
  1024 => x"c087c602",
  1025 => x"f105a9fb",
  1026 => x"26487187",
  1027 => x"5b5e0e4f",
  1028 => x"4b710e5c",
  1029 => x"f8fe4cc0",
  1030 => x"99497087",
  1031 => x"87f9c002",
  1032 => x"02a9ecc0",
  1033 => x"c087f2c0",
  1034 => x"c002a9fb",
  1035 => x"66cc87eb",
  1036 => x"c703acb7",
  1037 => x"0266d087",
  1038 => x"537187c2",
  1039 => x"c2029971",
  1040 => x"fe84c187",
  1041 => x"497087cb",
  1042 => x"87cd0299",
  1043 => x"02a9ecc0",
  1044 => x"fbc087c7",
  1045 => x"d5ff05a9",
  1046 => x"0266d087",
  1047 => x"97c087c3",
  1048 => x"a9ecc07b",
  1049 => x"7487c405",
  1050 => x"7487c54a",
  1051 => x"8a0ac04a",
  1052 => x"4c264872",
  1053 => x"4f264b26",
  1054 => x"87d5fd1e",
  1055 => x"f0c04970",
  1056 => x"87c904a9",
  1057 => x"01a9f9c0",
  1058 => x"f0c087c3",
  1059 => x"a9c1c189",
  1060 => x"c187c904",
  1061 => x"c301a9da",
  1062 => x"89f7c087",
  1063 => x"4f264871",
  1064 => x"5c5b5e0e",
  1065 => x"86f80e5d",
  1066 => x"7ec04c71",
  1067 => x"c087edfc",
  1068 => x"c0c5c14b",
  1069 => x"c049bf97",
  1070 => x"87cf04a9",
  1071 => x"c187fafc",
  1072 => x"c0c5c183",
  1073 => x"ab49bf97",
  1074 => x"c187f106",
  1075 => x"bf97c0c5",
  1076 => x"fb87cf02",
  1077 => x"497087fb",
  1078 => x"87c60299",
  1079 => x"05a9ecc0",
  1080 => x"4bc087f1",
  1081 => x"7087eafb",
  1082 => x"87e5fb4d",
  1083 => x"fb58a6c8",
  1084 => x"4a7087df",
  1085 => x"a4c883c1",
  1086 => x"49699749",
  1087 => x"87da05ad",
  1088 => x"9749a4c9",
  1089 => x"66c44969",
  1090 => x"87ce05a9",
  1091 => x"9749a4ca",
  1092 => x"05aa4969",
  1093 => x"7ec187c4",
  1094 => x"ecc087d0",
  1095 => x"87c602ad",
  1096 => x"05adfbc0",
  1097 => x"4bc087c4",
  1098 => x"026e7ec1",
  1099 => x"fa87f5fe",
  1100 => x"487387fe",
  1101 => x"4d268ef8",
  1102 => x"4b264c26",
  1103 => x"00004f26",
  1104 => x"1e731e00",
  1105 => x"c84bd4ff",
  1106 => x"d0ff4a66",
  1107 => x"78c5c848",
  1108 => x"c148d4ff",
  1109 => x"7b1178d4",
  1110 => x"f9058ac1",
  1111 => x"48d0ff87",
  1112 => x"4b2678c4",
  1113 => x"5e0e4f26",
  1114 => x"0e5d5c5b",
  1115 => x"7e7186f8",
  1116 => x"f7c21e6e",
  1117 => x"dfff49d4",
  1118 => x"86c487df",
  1119 => x"c4029870",
  1120 => x"f4c187e4",
  1121 => x"6e4cbfc8",
  1122 => x"87d4fc49",
  1123 => x"7058a6c8",
  1124 => x"87c50598",
  1125 => x"c148a6c4",
  1126 => x"48d0ff78",
  1127 => x"d4ff78c5",
  1128 => x"78d5c148",
  1129 => x"c14966c4",
  1130 => x"c131c689",
  1131 => x"bf97c0f4",
  1132 => x"b071484a",
  1133 => x"7808d4ff",
  1134 => x"c448d0ff",
  1135 => x"d0f7c278",
  1136 => x"d049bf97",
  1137 => x"87dd0299",
  1138 => x"d4ff78c5",
  1139 => x"78d6c148",
  1140 => x"d4ff4ac0",
  1141 => x"78ffc348",
  1142 => x"e0c082c1",
  1143 => x"87f204aa",
  1144 => x"c448d0ff",
  1145 => x"48d4ff78",
  1146 => x"ff78ffc3",
  1147 => x"78c548d0",
  1148 => x"c148d4ff",
  1149 => x"78c178d3",
  1150 => x"c448d0ff",
  1151 => x"acb7c078",
  1152 => x"87cbc206",
  1153 => x"bfdcf7c2",
  1154 => x"7e748c4b",
  1155 => x"c1029b73",
  1156 => x"c0c887dd",
  1157 => x"b7c08b4d",
  1158 => x"87c603ab",
  1159 => x"4da3c0c8",
  1160 => x"f7c24bc0",
  1161 => x"49bf97d0",
  1162 => x"cf0299d0",
  1163 => x"c21ec087",
  1164 => x"e249d4f7",
  1165 => x"86c487e1",
  1166 => x"87d84c70",
  1167 => x"1ed4eac2",
  1168 => x"49d4f7c2",
  1169 => x"7087d0e2",
  1170 => x"c21e754c",
  1171 => x"fb49d4ea",
  1172 => x"86c887ef",
  1173 => x"c5059c74",
  1174 => x"c148c087",
  1175 => x"1ec187ca",
  1176 => x"49d4f7c2",
  1177 => x"c487d5e0",
  1178 => x"059b7386",
  1179 => x"6e87e3fe",
  1180 => x"acb7c04c",
  1181 => x"c287d106",
  1182 => x"c048d4f7",
  1183 => x"c080d078",
  1184 => x"c280f478",
  1185 => x"78bfe0f7",
  1186 => x"01acb7c0",
  1187 => x"ff87f5fd",
  1188 => x"78c548d0",
  1189 => x"c148d4ff",
  1190 => x"78c078d3",
  1191 => x"c448d0ff",
  1192 => x"c048c178",
  1193 => x"48c087c2",
  1194 => x"4d268ef8",
  1195 => x"4b264c26",
  1196 => x"5e0e4f26",
  1197 => x"0e5d5c5b",
  1198 => x"4d7186fc",
  1199 => x"ad4c4bc0",
  1200 => x"87e8c004",
  1201 => x"1ee0c2c1",
  1202 => x"c4029c74",
  1203 => x"c24ac087",
  1204 => x"724ac187",
  1205 => x"87e0eb49",
  1206 => x"7e7086c4",
  1207 => x"056e83c1",
  1208 => x"4b7587c2",
  1209 => x"ab7584c1",
  1210 => x"87d8ff06",
  1211 => x"8efc486e",
  1212 => x"4c264d26",
  1213 => x"4f264b26",
  1214 => x"5c5b5e0e",
  1215 => x"cc4b710e",
  1216 => x"87d80266",
  1217 => x"8cf0c04c",
  1218 => x"7487d802",
  1219 => x"028ac14a",
  1220 => x"028a87d1",
  1221 => x"028a87cd",
  1222 => x"87d987c9",
  1223 => x"c5f94973",
  1224 => x"7487d287",
  1225 => x"c149c01e",
  1226 => x"7487fdd9",
  1227 => x"c149731e",
  1228 => x"c887f5d9",
  1229 => x"264c2686",
  1230 => x"0e4f264b",
  1231 => x"5d5c5b5e",
  1232 => x"7186fc0e",
  1233 => x"91de494c",
  1234 => x"4df4f8c2",
  1235 => x"6d978571",
  1236 => x"87dcc102",
  1237 => x"bfe4f8c2",
  1238 => x"71817449",
  1239 => x"7087d3fd",
  1240 => x"0298487e",
  1241 => x"c287f2c0",
  1242 => x"704be8f8",
  1243 => x"fe49cb4a",
  1244 => x"7487f1f6",
  1245 => x"c193cc4b",
  1246 => x"c483ccf4",
  1247 => x"fccec183",
  1248 => x"c149747b",
  1249 => x"7587e9c4",
  1250 => x"c4f4c17b",
  1251 => x"1e49bf97",
  1252 => x"49e8f8c2",
  1253 => x"c487e1fd",
  1254 => x"c1497486",
  1255 => x"c087d1c4",
  1256 => x"ecc5c149",
  1257 => x"ccf7c287",
  1258 => x"4950c048",
  1259 => x"87cbe2c0",
  1260 => x"4d268efc",
  1261 => x"4b264c26",
  1262 => x"00004f26",
  1263 => x"64616f4c",
  1264 => x"2e676e69",
  1265 => x"1e002e2e",
  1266 => x"4b711e73",
  1267 => x"e4f8c249",
  1268 => x"fb7181bf",
  1269 => x"4a7087dc",
  1270 => x"87c4029a",
  1271 => x"87dee649",
  1272 => x"48e4f8c2",
  1273 => x"497378c0",
  1274 => x"2687fac1",
  1275 => x"1e4f264b",
  1276 => x"4b711e73",
  1277 => x"024aa3c4",
  1278 => x"c187d0c1",
  1279 => x"87dc028a",
  1280 => x"f2c0028a",
  1281 => x"c1058a87",
  1282 => x"f8c287d3",
  1283 => x"c102bfe4",
  1284 => x"c14887cb",
  1285 => x"e8f8c288",
  1286 => x"87c1c158",
  1287 => x"bfe4f8c2",
  1288 => x"c289c649",
  1289 => x"c059e8f8",
  1290 => x"c003a9b7",
  1291 => x"f8c287ef",
  1292 => x"78c048e4",
  1293 => x"c287e6c0",
  1294 => x"02bfe0f8",
  1295 => x"f8c287df",
  1296 => x"c148bfe4",
  1297 => x"e8f8c280",
  1298 => x"c287d258",
  1299 => x"02bfe0f8",
  1300 => x"f8c287cb",
  1301 => x"c648bfe4",
  1302 => x"e8f8c280",
  1303 => x"c4497358",
  1304 => x"264b2687",
  1305 => x"5b5e0e4f",
  1306 => x"f00e5d5c",
  1307 => x"59a6d086",
  1308 => x"4dd4eac2",
  1309 => x"f8c24cc0",
  1310 => x"78c148e0",
  1311 => x"c048a6c8",
  1312 => x"c27e7578",
  1313 => x"48bfe4f8",
  1314 => x"c106a8c0",
  1315 => x"a6c887c0",
  1316 => x"c27e755c",
  1317 => x"9848d4ea",
  1318 => x"87f2c002",
  1319 => x"c14d66c4",
  1320 => x"cc1ee0c2",
  1321 => x"87c40266",
  1322 => x"87c24cc0",
  1323 => x"49744cc1",
  1324 => x"c487c5e4",
  1325 => x"c17e7086",
  1326 => x"4866c885",
  1327 => x"a6cc80c1",
  1328 => x"e4f8c258",
  1329 => x"c503adbf",
  1330 => x"ff056e87",
  1331 => x"4d6e87d1",
  1332 => x"9d754cc0",
  1333 => x"87dcc302",
  1334 => x"1ee0c2c1",
  1335 => x"c70266cc",
  1336 => x"48a6c887",
  1337 => x"87c578c0",
  1338 => x"c148a6c8",
  1339 => x"4966c878",
  1340 => x"c487c5e3",
  1341 => x"487e7086",
  1342 => x"e4c20298",
  1343 => x"81cb4987",
  1344 => x"d0496997",
  1345 => x"d4c10299",
  1346 => x"cc497487",
  1347 => x"ccf4c191",
  1348 => x"c7cfc181",
  1349 => x"c381c879",
  1350 => x"497451ff",
  1351 => x"f8c291de",
  1352 => x"85714df4",
  1353 => x"7d97c1c2",
  1354 => x"c049a5c1",
  1355 => x"f2c251e0",
  1356 => x"02bf97e4",
  1357 => x"84c187d2",
  1358 => x"c24ba5c2",
  1359 => x"db4ae4f2",
  1360 => x"dfeffe49",
  1361 => x"87d9c187",
  1362 => x"c049a5cd",
  1363 => x"c284c151",
  1364 => x"4a6e4ba5",
  1365 => x"effe49cb",
  1366 => x"c4c187ca",
  1367 => x"cc497487",
  1368 => x"ccf4c191",
  1369 => x"fbccc181",
  1370 => x"e4f2c279",
  1371 => x"d802bf97",
  1372 => x"de497487",
  1373 => x"c284c191",
  1374 => x"714bf4f8",
  1375 => x"e4f2c283",
  1376 => x"fe49dd4a",
  1377 => x"d887ddee",
  1378 => x"de4b7487",
  1379 => x"f4f8c293",
  1380 => x"49a3cb83",
  1381 => x"84c151c0",
  1382 => x"cb4a6e73",
  1383 => x"c3eefe49",
  1384 => x"4866c887",
  1385 => x"a6cc80c1",
  1386 => x"03acc758",
  1387 => x"6e87c5c0",
  1388 => x"87e4fc05",
  1389 => x"c003acc7",
  1390 => x"f8c287e4",
  1391 => x"78c048e0",
  1392 => x"91cc4974",
  1393 => x"81ccf4c1",
  1394 => x"79fbccc1",
  1395 => x"91de4974",
  1396 => x"81f4f8c2",
  1397 => x"84c151c0",
  1398 => x"ff04acc7",
  1399 => x"f5c187dc",
  1400 => x"50c048e8",
  1401 => x"d9c180f7",
  1402 => x"d8c140d5",
  1403 => x"80c878c8",
  1404 => x"78efcfc1",
  1405 => x"c04966cc",
  1406 => x"f087f5fa",
  1407 => x"264d268e",
  1408 => x"264b264c",
  1409 => x"0000004f",
  1410 => x"61422080",
  1411 => x"1e006b63",
  1412 => x"4b711e73",
  1413 => x"c191cc49",
  1414 => x"c881ccf4",
  1415 => x"f4c14aa1",
  1416 => x"501248c0",
  1417 => x"c14aa1c9",
  1418 => x"1248c0c5",
  1419 => x"c181ca50",
  1420 => x"1148c4f4",
  1421 => x"c4f4c150",
  1422 => x"1e49bf97",
  1423 => x"f7f249c0",
  1424 => x"f8497387",
  1425 => x"8efc87df",
  1426 => x"4f264b26",
  1427 => x"c049c01e",
  1428 => x"2687fefa",
  1429 => x"4a711e4f",
  1430 => x"c191cc49",
  1431 => x"c881ccf4",
  1432 => x"ccf7c281",
  1433 => x"c0501148",
  1434 => x"fe49a2f0",
  1435 => x"c087dde8",
  1436 => x"87c7d749",
  1437 => x"ff1e4f26",
  1438 => x"ffc34ad4",
  1439 => x"48d0ff7a",
  1440 => x"de78e1c0",
  1441 => x"487a717a",
  1442 => x"7028b7c8",
  1443 => x"d048717a",
  1444 => x"7a7028b7",
  1445 => x"b7d84871",
  1446 => x"ff7a7028",
  1447 => x"e0c048d0",
  1448 => x"0e4f2678",
  1449 => x"5d5c5b5e",
  1450 => x"7186f40e",
  1451 => x"91cc494d",
  1452 => x"81ccf4c1",
  1453 => x"ca4aa1c8",
  1454 => x"a6c47ea1",
  1455 => x"c8f7c248",
  1456 => x"976e78bf",
  1457 => x"66c44bbf",
  1458 => x"122c734c",
  1459 => x"58a6cc48",
  1460 => x"84c19c70",
  1461 => x"699781c9",
  1462 => x"04acb749",
  1463 => x"4cc087c2",
  1464 => x"4abf976e",
  1465 => x"724966c8",
  1466 => x"c4b9ff31",
  1467 => x"48749966",
  1468 => x"4a703072",
  1469 => x"ccf7c2b1",
  1470 => x"f9fd7159",
  1471 => x"c21ec787",
  1472 => x"1ebfdcf8",
  1473 => x"1eccf4c1",
  1474 => x"97ccf7c2",
  1475 => x"f4c149bf",
  1476 => x"c0497587",
  1477 => x"e887d9f6",
  1478 => x"264d268e",
  1479 => x"264b264c",
  1480 => x"1e731e4f",
  1481 => x"fd494b71",
  1482 => x"497387f9",
  1483 => x"2687f4fd",
  1484 => x"1e4f264b",
  1485 => x"4b711e73",
  1486 => x"024aa3c2",
  1487 => x"8ac187d6",
  1488 => x"87e2c005",
  1489 => x"bfdcf8c2",
  1490 => x"4887db02",
  1491 => x"f8c288c1",
  1492 => x"87d258e0",
  1493 => x"bfe0f8c2",
  1494 => x"c287cb02",
  1495 => x"48bfdcf8",
  1496 => x"f8c280c1",
  1497 => x"1ec758e0",
  1498 => x"bfdcf8c2",
  1499 => x"ccf4c11e",
  1500 => x"ccf7c21e",
  1501 => x"cc49bf97",
  1502 => x"c0497387",
  1503 => x"f487f1f4",
  1504 => x"264b268e",
  1505 => x"5b5e0e4f",
  1506 => x"ff0e5d5c",
  1507 => x"e4c086cc",
  1508 => x"a6cc59a6",
  1509 => x"c478c048",
  1510 => x"c478c080",
  1511 => x"66c8c180",
  1512 => x"c180c478",
  1513 => x"c180c478",
  1514 => x"e0f8c278",
  1515 => x"e078c148",
  1516 => x"c4e187ea",
  1517 => x"87d9e087",
  1518 => x"fbc04c70",
  1519 => x"f3c102ac",
  1520 => x"66e0c087",
  1521 => x"87e8c105",
  1522 => x"4a66c4c1",
  1523 => x"7e6a82c4",
  1524 => x"48dcf0c1",
  1525 => x"4120496e",
  1526 => x"51104120",
  1527 => x"4866c4c1",
  1528 => x"78cfd8c1",
  1529 => x"81c7496a",
  1530 => x"c4c15174",
  1531 => x"81c84966",
  1532 => x"a6d851c1",
  1533 => x"c178c248",
  1534 => x"c94966c4",
  1535 => x"c151c081",
  1536 => x"ca4966c4",
  1537 => x"c151c081",
  1538 => x"6a1ed81e",
  1539 => x"ff81c849",
  1540 => x"c887fadf",
  1541 => x"66c8c186",
  1542 => x"01a8c048",
  1543 => x"a6d087c7",
  1544 => x"cf78c148",
  1545 => x"66c8c187",
  1546 => x"d888c148",
  1547 => x"87c458a6",
  1548 => x"87c5dfff",
  1549 => x"cd029c74",
  1550 => x"66d087d9",
  1551 => x"66ccc148",
  1552 => x"cecd03a8",
  1553 => x"48a6c887",
  1554 => x"ff7e78c0",
  1555 => x"7087c2de",
  1556 => x"acd0c14c",
  1557 => x"87e7c205",
  1558 => x"6e48a6c4",
  1559 => x"87d8e078",
  1560 => x"cc487e70",
  1561 => x"c506a866",
  1562 => x"48a6cc87",
  1563 => x"ddff786e",
  1564 => x"4c7087df",
  1565 => x"05acecc0",
  1566 => x"d087eec1",
  1567 => x"91cc4966",
  1568 => x"8166c4c1",
  1569 => x"6a4aa1c4",
  1570 => x"4aa1c84d",
  1571 => x"d9c1526e",
  1572 => x"dcff79d5",
  1573 => x"4c7087fb",
  1574 => x"87d9029c",
  1575 => x"02acfbc0",
  1576 => x"557487d3",
  1577 => x"87e9dcff",
  1578 => x"029c4c70",
  1579 => x"fbc087c7",
  1580 => x"edff05ac",
  1581 => x"55e0c087",
  1582 => x"c055c1c2",
  1583 => x"e0c07d97",
  1584 => x"66c44866",
  1585 => x"87db05a8",
  1586 => x"d44866d0",
  1587 => x"ca04a866",
  1588 => x"4866d087",
  1589 => x"a6d480c1",
  1590 => x"d487c858",
  1591 => x"88c14866",
  1592 => x"ff58a6d8",
  1593 => x"7087eadb",
  1594 => x"acd0c14c",
  1595 => x"dc87c905",
  1596 => x"80c14866",
  1597 => x"58a6e0c0",
  1598 => x"02acd0c1",
  1599 => x"6e87d9fd",
  1600 => x"66e0c048",
  1601 => x"eac905a8",
  1602 => x"a6e4c087",
  1603 => x"7478c048",
  1604 => x"88fbc048",
  1605 => x"7058a6c8",
  1606 => x"dcc90298",
  1607 => x"88cb4887",
  1608 => x"7058a6c8",
  1609 => x"cec10298",
  1610 => x"88c94887",
  1611 => x"7058a6c8",
  1612 => x"fec30298",
  1613 => x"88c44887",
  1614 => x"7058a6c8",
  1615 => x"87cf0298",
  1616 => x"c888c148",
  1617 => x"987058a6",
  1618 => x"87e7c302",
  1619 => x"c887dbc8",
  1620 => x"f0c048a6",
  1621 => x"f8d9ff78",
  1622 => x"c04c7087",
  1623 => x"c302acec",
  1624 => x"5ca6cc87",
  1625 => x"02acecc0",
  1626 => x"d9ff87cd",
  1627 => x"4c7087e3",
  1628 => x"05acecc0",
  1629 => x"c087f3ff",
  1630 => x"c002acec",
  1631 => x"d9ff87c4",
  1632 => x"1ec087cf",
  1633 => x"66d81eca",
  1634 => x"c191cc49",
  1635 => x"714866cc",
  1636 => x"58a6cc80",
  1637 => x"c44866c8",
  1638 => x"58a6d080",
  1639 => x"49bf66cc",
  1640 => x"87e9d9ff",
  1641 => x"1ede1ec1",
  1642 => x"49bf66d4",
  1643 => x"87ddd9ff",
  1644 => x"497086d0",
  1645 => x"8808c048",
  1646 => x"58a6ecc0",
  1647 => x"c006a8c0",
  1648 => x"e8c087ee",
  1649 => x"a8dd4866",
  1650 => x"87e4c003",
  1651 => x"49bf66c4",
  1652 => x"8166e8c0",
  1653 => x"c051e0c0",
  1654 => x"c14966e8",
  1655 => x"bf66c481",
  1656 => x"51c1c281",
  1657 => x"4966e8c0",
  1658 => x"66c481c2",
  1659 => x"51c081bf",
  1660 => x"d8c1486e",
  1661 => x"496e78cf",
  1662 => x"66d881c8",
  1663 => x"c9496e51",
  1664 => x"5166dc81",
  1665 => x"81ca496e",
  1666 => x"d85166c8",
  1667 => x"80c14866",
  1668 => x"d058a6dc",
  1669 => x"66d44866",
  1670 => x"cbc004a8",
  1671 => x"4866d087",
  1672 => x"a6d480c1",
  1673 => x"87d1c558",
  1674 => x"c14866d4",
  1675 => x"58a6d888",
  1676 => x"ff87c6c5",
  1677 => x"c087c1d9",
  1678 => x"ff58a6ec",
  1679 => x"c087f9d8",
  1680 => x"c058a6f0",
  1681 => x"c005a8ec",
  1682 => x"48a687c9",
  1683 => x"7866e8c0",
  1684 => x"ff87c4c0",
  1685 => x"d087fad5",
  1686 => x"91cc4966",
  1687 => x"4866c4c1",
  1688 => x"a6c88071",
  1689 => x"4a66c458",
  1690 => x"66c482c8",
  1691 => x"c081ca49",
  1692 => x"c05166e8",
  1693 => x"c14966ec",
  1694 => x"66e8c081",
  1695 => x"7148c189",
  1696 => x"c1497030",
  1697 => x"7a977189",
  1698 => x"bfc8f7c2",
  1699 => x"66e8c049",
  1700 => x"4a6a9729",
  1701 => x"c0987148",
  1702 => x"c458a6f4",
  1703 => x"80c44866",
  1704 => x"c858a6cc",
  1705 => x"c04dbf66",
  1706 => x"6e4866e0",
  1707 => x"c5c002a8",
  1708 => x"c07ec087",
  1709 => x"7ec187c2",
  1710 => x"e0c01e6e",
  1711 => x"ff49751e",
  1712 => x"c887cad5",
  1713 => x"c04c7086",
  1714 => x"c106acb7",
  1715 => x"857487d4",
  1716 => x"49bf66c8",
  1717 => x"7581e0c0",
  1718 => x"f0c14b89",
  1719 => x"fe714ae8",
  1720 => x"c287c1d9",
  1721 => x"c07e7585",
  1722 => x"c14866e4",
  1723 => x"a6e8c080",
  1724 => x"66f0c058",
  1725 => x"7081c149",
  1726 => x"c5c002a9",
  1727 => x"c04dc087",
  1728 => x"4dc187c2",
  1729 => x"66cc1e75",
  1730 => x"e0c049bf",
  1731 => x"8966c481",
  1732 => x"66c81e71",
  1733 => x"f4d3ff49",
  1734 => x"c086c887",
  1735 => x"ff01a8b7",
  1736 => x"e4c087c5",
  1737 => x"d3c00266",
  1738 => x"4966c487",
  1739 => x"e4c081c9",
  1740 => x"66c45166",
  1741 => x"e3dac148",
  1742 => x"87cec078",
  1743 => x"c94966c4",
  1744 => x"c451c281",
  1745 => x"dcc14866",
  1746 => x"66d078e1",
  1747 => x"a866d448",
  1748 => x"87cbc004",
  1749 => x"c14866d0",
  1750 => x"58a6d480",
  1751 => x"d487dac0",
  1752 => x"88c14866",
  1753 => x"c058a6d8",
  1754 => x"d2ff87cf",
  1755 => x"4c7087cb",
  1756 => x"ff87c6c0",
  1757 => x"7087c2d2",
  1758 => x"4866dc4c",
  1759 => x"e0c080c1",
  1760 => x"9c7458a6",
  1761 => x"87cbc002",
  1762 => x"c14866d0",
  1763 => x"04a866cc",
  1764 => x"d087f2f2",
  1765 => x"a8c74866",
  1766 => x"87e1c003",
  1767 => x"c24c66d0",
  1768 => x"c048e0f8",
  1769 => x"cc497478",
  1770 => x"66c4c191",
  1771 => x"4aa1c481",
  1772 => x"52c04a6a",
  1773 => x"c784c179",
  1774 => x"e2ff04ac",
  1775 => x"66e0c087",
  1776 => x"87e2c002",
  1777 => x"4966c4c1",
  1778 => x"c181d4c1",
  1779 => x"c14a66c4",
  1780 => x"52c082dc",
  1781 => x"79d5d9c1",
  1782 => x"4966c4c1",
  1783 => x"c181d8c1",
  1784 => x"c079ecf0",
  1785 => x"c4c187d6",
  1786 => x"d4c14966",
  1787 => x"66c4c181",
  1788 => x"82d8c14a",
  1789 => x"7af4f0c1",
  1790 => x"79ccd9c1",
  1791 => x"4966c4c1",
  1792 => x"c181e0c1",
  1793 => x"ff79f3dc",
  1794 => x"cc87e5cf",
  1795 => x"ccff4866",
  1796 => x"264d268e",
  1797 => x"264b264c",
  1798 => x"0000004f",
  1799 => x"64616f4c",
  1800 => x"202e2a20",
  1801 => x"00000000",
  1802 => x"0000203a",
  1803 => x"61422080",
  1804 => x"00006b63",
  1805 => x"78452080",
  1806 => x"1e007469",
  1807 => x"f8c21ec7",
  1808 => x"c11ebfdc",
  1809 => x"c21eccf4",
  1810 => x"bf97ccf7",
  1811 => x"87f5ec49",
  1812 => x"49ccf4c1",
  1813 => x"87e6e2c0",
  1814 => x"4f268ef4",
  1815 => x"c81e731e",
  1816 => x"f5c187c3",
  1817 => x"f3c148e4",
  1818 => x"e8fe78ec",
  1819 => x"e2c049a0",
  1820 => x"49c787cc",
  1821 => x"87f8e0c0",
  1822 => x"e2c049c1",
  1823 => x"d4ff87d3",
  1824 => x"78ffc348",
  1825 => x"48e8f8c2",
  1826 => x"ddfe50c0",
  1827 => x"987087e2",
  1828 => x"fe87cd02",
  1829 => x"7087dee7",
  1830 => x"87c40298",
  1831 => x"87c24ac1",
  1832 => x"9a724ac0",
  1833 => x"c187c802",
  1834 => x"fe49f8f3",
  1835 => x"c287f8cf",
  1836 => x"c048dcf8",
  1837 => x"ccf7c278",
  1838 => x"4950c048",
  1839 => x"c087fcfd",
  1840 => x"7087eaf5",
  1841 => x"cb029b4b",
  1842 => x"e8f5c187",
  1843 => x"df49c75b",
  1844 => x"87c687de",
  1845 => x"e0c049c0",
  1846 => x"c2c387f7",
  1847 => x"d8e2c087",
  1848 => x"ecefc087",
  1849 => x"87f5ff87",
  1850 => x"4f264b26",
  1851 => x"746f6f42",
  1852 => x"2e676e69",
  1853 => x"00002e2e",
  1854 => x"4f204453",
  1855 => x"0000004b",
  1856 => x"00000000",
  1857 => x"00000000",
  1858 => x"00000001",
  1859 => x"0000133b",
  1860 => x"00002e34",
  1861 => x"00000000",
  1862 => x"0000133b",
  1863 => x"00002e52",
  1864 => x"00000000",
  1865 => x"0000133b",
  1866 => x"00002e70",
  1867 => x"00000000",
  1868 => x"0000133b",
  1869 => x"00002e8e",
  1870 => x"00000000",
  1871 => x"0000133b",
  1872 => x"00002eac",
  1873 => x"00000000",
  1874 => x"0000133b",
  1875 => x"00002eca",
  1876 => x"00000000",
  1877 => x"0000133b",
  1878 => x"00002ee8",
  1879 => x"00000000",
  1880 => x"00001655",
  1881 => x"00000000",
  1882 => x"00000000",
  1883 => x"000013ef",
  1884 => x"00000000",
  1885 => x"00000000",
  1886 => x"db86fc1e",
  1887 => x"fc7e7087",
  1888 => x"1e4f268e",
  1889 => x"c048f0fe",
  1890 => x"7909cd78",
  1891 => x"1e4f2609",
  1892 => x"49f8f5c1",
  1893 => x"4f2687ed",
  1894 => x"bff0fe1e",
  1895 => x"1e4f2648",
  1896 => x"c148f0fe",
  1897 => x"1e4f2678",
  1898 => x"c048f0fe",
  1899 => x"1e4f2678",
  1900 => x"52c04a71",
  1901 => x"0e4f2651",
  1902 => x"5d5c5b5e",
  1903 => x"7186f40e",
  1904 => x"7e6d974d",
  1905 => x"974ca5c1",
  1906 => x"a6c8486c",
  1907 => x"c4486e58",
  1908 => x"c505a866",
  1909 => x"c048ff87",
  1910 => x"caff87e6",
  1911 => x"49a5c287",
  1912 => x"714b6c97",
  1913 => x"6b974ba3",
  1914 => x"7e6c974b",
  1915 => x"80c1486e",
  1916 => x"c758a6c8",
  1917 => x"58a6cc98",
  1918 => x"fe7c9770",
  1919 => x"487387e1",
  1920 => x"4d268ef4",
  1921 => x"4b264c26",
  1922 => x"5e0e4f26",
  1923 => x"f40e5c5b",
  1924 => x"d84c7186",
  1925 => x"ffc34a66",
  1926 => x"4ba4c29a",
  1927 => x"73496c97",
  1928 => x"517249a1",
  1929 => x"6e7e6c97",
  1930 => x"c880c148",
  1931 => x"98c758a6",
  1932 => x"7058a6cc",
  1933 => x"268ef454",
  1934 => x"264b264c",
  1935 => x"86fc1e4f",
  1936 => x"e087e4fd",
  1937 => x"c0494abf",
  1938 => x"0299c0e0",
  1939 => x"1e7287cb",
  1940 => x"49c8fcc2",
  1941 => x"c487f3fe",
  1942 => x"87fcfc86",
  1943 => x"fefc7e70",
  1944 => x"268efc87",
  1945 => x"fcc21e4f",
  1946 => x"c2fd49c8",
  1947 => x"fdf8c187",
  1948 => x"87cffc49",
  1949 => x"2687edc3",
  1950 => x"5b5e0e4f",
  1951 => x"fc0e5d5c",
  1952 => x"ff7e7186",
  1953 => x"fcc24dd4",
  1954 => x"eafc49c8",
  1955 => x"c04b7087",
  1956 => x"c204abb7",
  1957 => x"f0c387f8",
  1958 => x"87c905ab",
  1959 => x"48dcfdc1",
  1960 => x"d9c278c1",
  1961 => x"abe0c387",
  1962 => x"c187c905",
  1963 => x"c148e0fd",
  1964 => x"87cac278",
  1965 => x"bfe0fdc1",
  1966 => x"c287c602",
  1967 => x"c24ca3c0",
  1968 => x"c14c7387",
  1969 => x"02bfdcfd",
  1970 => x"7487e0c0",
  1971 => x"29b7c449",
  1972 => x"f8fec191",
  1973 => x"cf4a7481",
  1974 => x"c192c29a",
  1975 => x"70307248",
  1976 => x"72baff4a",
  1977 => x"70986948",
  1978 => x"7487db79",
  1979 => x"29b7c449",
  1980 => x"f8fec191",
  1981 => x"cf4a7481",
  1982 => x"c392c29a",
  1983 => x"70307248",
  1984 => x"b069484a",
  1985 => x"056e7970",
  1986 => x"ff87e7c0",
  1987 => x"e1c848d0",
  1988 => x"c17dc578",
  1989 => x"02bfe0fd",
  1990 => x"e0c387c3",
  1991 => x"dcfdc17d",
  1992 => x"87c302bf",
  1993 => x"737df0c3",
  1994 => x"48d0ff7d",
  1995 => x"c078e1c8",
  1996 => x"fdc178e0",
  1997 => x"78c048e0",
  1998 => x"48dcfdc1",
  1999 => x"fcc278c0",
  2000 => x"f2f949c8",
  2001 => x"c04b7087",
  2002 => x"fd03abb7",
  2003 => x"48c087c8",
  2004 => x"4d268efc",
  2005 => x"4b264c26",
  2006 => x"00004f26",
  2007 => x"00000000",
  2008 => x"00000000",
  2009 => x"724ac01e",
  2010 => x"c191c449",
  2011 => x"c081f8fe",
  2012 => x"d082c179",
  2013 => x"ee04aab7",
  2014 => x"0e4f2687",
  2015 => x"5d5c5b5e",
  2016 => x"f84d710e",
  2017 => x"4a7587e1",
  2018 => x"922ab7c4",
  2019 => x"82f8fec1",
  2020 => x"9ccf4c75",
  2021 => x"496a94c2",
  2022 => x"c32b744b",
  2023 => x"7448c29b",
  2024 => x"ff4c7030",
  2025 => x"714874bc",
  2026 => x"f77a7098",
  2027 => x"487387f1",
  2028 => x"4c264d26",
  2029 => x"4f264b26",
  2030 => x"00000000",
  2031 => x"00000000",
  2032 => x"00000000",
  2033 => x"00000000",
  2034 => x"00000000",
  2035 => x"00000000",
  2036 => x"00000000",
  2037 => x"00000000",
  2038 => x"00000000",
  2039 => x"00000000",
  2040 => x"00000000",
  2041 => x"00000000",
  2042 => x"00000000",
  2043 => x"00000000",
  2044 => x"00000000",
  2045 => x"00000000",
  2046 => x"48d0ff1e",
  2047 => x"7178e1c8",
  2048 => x"08d4ff48",
  2049 => x"1e4f2678",
  2050 => x"c848d0ff",
  2051 => x"487178e1",
  2052 => x"7808d4ff",
  2053 => x"ff4866c4",
  2054 => x"267808d4",
  2055 => x"4a711e4f",
  2056 => x"1e4966c4",
  2057 => x"deff4972",
  2058 => x"48d0ff87",
  2059 => x"fc78e0c0",
  2060 => x"1e4f268e",
  2061 => x"4a711e73",
  2062 => x"abb7c24b",
  2063 => x"a387c803",
  2064 => x"ffc34a49",
  2065 => x"ce87c79a",
  2066 => x"c34a49a3",
  2067 => x"66c89aff",
  2068 => x"49721e49",
  2069 => x"fc87c6ff",
  2070 => x"264b268e",
  2071 => x"d0ff1e4f",
  2072 => x"78c9c848",
  2073 => x"d4ff4871",
  2074 => x"4f267808",
  2075 => x"494a711e",
  2076 => x"d0ff87eb",
  2077 => x"2678c848",
  2078 => x"1e731e4f",
  2079 => x"fcc24b71",
  2080 => x"c302bfe0",
  2081 => x"87ebc287",
  2082 => x"c848d0ff",
  2083 => x"487378c9",
  2084 => x"ffb0e0c0",
  2085 => x"c27808d4",
  2086 => x"c048d4fc",
  2087 => x"0266c878",
  2088 => x"ffc387c5",
  2089 => x"c087c249",
  2090 => x"dcfcc249",
  2091 => x"0266cc59",
  2092 => x"d5c587c6",
  2093 => x"87c44ad5",
  2094 => x"4affffcf",
  2095 => x"5ae0fcc2",
  2096 => x"48e0fcc2",
  2097 => x"4b2678c1",
  2098 => x"5e0e4f26",
  2099 => x"0e5d5c5b",
  2100 => x"fcc24d71",
  2101 => x"754bbfdc",
  2102 => x"87cb029d",
  2103 => x"c291c849",
  2104 => x"714af0c1",
  2105 => x"c287c482",
  2106 => x"c04af0c5",
  2107 => x"7349124c",
  2108 => x"d8fcc299",
  2109 => x"b87148bf",
  2110 => x"7808d4ff",
  2111 => x"842bb7c1",
  2112 => x"04acb7c8",
  2113 => x"fcc287e7",
  2114 => x"c848bfd4",
  2115 => x"d8fcc280",
  2116 => x"264d2658",
  2117 => x"264b264c",
  2118 => x"1e731e4f",
  2119 => x"4a134b71",
  2120 => x"87cb029a",
  2121 => x"e1fe4972",
  2122 => x"9a4a1387",
  2123 => x"2687f505",
  2124 => x"1e4f264b",
  2125 => x"bfd4fcc2",
  2126 => x"d4fcc249",
  2127 => x"78a1c148",
  2128 => x"a9b7c0c4",
  2129 => x"ff87db03",
  2130 => x"fcc248d4",
  2131 => x"c278bfd8",
  2132 => x"49bfd4fc",
  2133 => x"48d4fcc2",
  2134 => x"c478a1c1",
  2135 => x"04a9b7c0",
  2136 => x"d0ff87e5",
  2137 => x"c278c848",
  2138 => x"c048e0fc",
  2139 => x"004f2678",
  2140 => x"00000000",
  2141 => x"00000000",
  2142 => x"5f000000",
  2143 => x"0000005f",
  2144 => x"00030300",
  2145 => x"00000303",
  2146 => x"147f7f14",
  2147 => x"00147f7f",
  2148 => x"6b2e2400",
  2149 => x"00123a6b",
  2150 => x"18366a4c",
  2151 => x"0032566c",
  2152 => x"594f7e30",
  2153 => x"40683a77",
  2154 => x"07040000",
  2155 => x"00000003",
  2156 => x"3e1c0000",
  2157 => x"00004163",
  2158 => x"63410000",
  2159 => x"00001c3e",
  2160 => x"1c3e2a08",
  2161 => x"082a3e1c",
  2162 => x"3e080800",
  2163 => x"0008083e",
  2164 => x"e0800000",
  2165 => x"00000060",
  2166 => x"08080800",
  2167 => x"00080808",
  2168 => x"60000000",
  2169 => x"00000060",
  2170 => x"18306040",
  2171 => x"0103060c",
  2172 => x"597f3e00",
  2173 => x"003e7f4d",
  2174 => x"7f060400",
  2175 => x"0000007f",
  2176 => x"71634200",
  2177 => x"00464f59",
  2178 => x"49632200",
  2179 => x"00367f49",
  2180 => x"13161c18",
  2181 => x"00107f7f",
  2182 => x"45672700",
  2183 => x"00397d45",
  2184 => x"4b7e3c00",
  2185 => x"00307949",
  2186 => x"71010100",
  2187 => x"00070f79",
  2188 => x"497f3600",
  2189 => x"00367f49",
  2190 => x"494f0600",
  2191 => x"001e3f69",
  2192 => x"66000000",
  2193 => x"00000066",
  2194 => x"e6800000",
  2195 => x"00000066",
  2196 => x"14080800",
  2197 => x"00222214",
  2198 => x"14141400",
  2199 => x"00141414",
  2200 => x"14222200",
  2201 => x"00080814",
  2202 => x"51030200",
  2203 => x"00060f59",
  2204 => x"5d417f3e",
  2205 => x"001e1f55",
  2206 => x"097f7e00",
  2207 => x"007e7f09",
  2208 => x"497f7f00",
  2209 => x"00367f49",
  2210 => x"633e1c00",
  2211 => x"00414141",
  2212 => x"417f7f00",
  2213 => x"001c3e63",
  2214 => x"497f7f00",
  2215 => x"00414149",
  2216 => x"097f7f00",
  2217 => x"00010109",
  2218 => x"417f3e00",
  2219 => x"007a7b49",
  2220 => x"087f7f00",
  2221 => x"007f7f08",
  2222 => x"7f410000",
  2223 => x"0000417f",
  2224 => x"40602000",
  2225 => x"003f7f40",
  2226 => x"1c087f7f",
  2227 => x"00416336",
  2228 => x"407f7f00",
  2229 => x"00404040",
  2230 => x"0c067f7f",
  2231 => x"007f7f06",
  2232 => x"0c067f7f",
  2233 => x"007f7f18",
  2234 => x"417f3e00",
  2235 => x"003e7f41",
  2236 => x"097f7f00",
  2237 => x"00060f09",
  2238 => x"61417f3e",
  2239 => x"00407e7f",
  2240 => x"097f7f00",
  2241 => x"00667f19",
  2242 => x"4d6f2600",
  2243 => x"00327b59",
  2244 => x"7f010100",
  2245 => x"0001017f",
  2246 => x"407f3f00",
  2247 => x"003f7f40",
  2248 => x"703f0f00",
  2249 => x"000f3f70",
  2250 => x"18307f7f",
  2251 => x"007f7f30",
  2252 => x"1c366341",
  2253 => x"4163361c",
  2254 => x"7c060301",
  2255 => x"0103067c",
  2256 => x"4d597161",
  2257 => x"00414347",
  2258 => x"7f7f0000",
  2259 => x"00004141",
  2260 => x"0c060301",
  2261 => x"40603018",
  2262 => x"41410000",
  2263 => x"00007f7f",
  2264 => x"03060c08",
  2265 => x"00080c06",
  2266 => x"80808080",
  2267 => x"00808080",
  2268 => x"03000000",
  2269 => x"00000407",
  2270 => x"54742000",
  2271 => x"00787c54",
  2272 => x"447f7f00",
  2273 => x"00387c44",
  2274 => x"447c3800",
  2275 => x"00004444",
  2276 => x"447c3800",
  2277 => x"007f7f44",
  2278 => x"547c3800",
  2279 => x"00185c54",
  2280 => x"7f7e0400",
  2281 => x"00000505",
  2282 => x"a4bc1800",
  2283 => x"007cfca4",
  2284 => x"047f7f00",
  2285 => x"00787c04",
  2286 => x"3d000000",
  2287 => x"0000407d",
  2288 => x"80808000",
  2289 => x"00007dfd",
  2290 => x"107f7f00",
  2291 => x"00446c38",
  2292 => x"3f000000",
  2293 => x"0000407f",
  2294 => x"180c7c7c",
  2295 => x"00787c0c",
  2296 => x"047c7c00",
  2297 => x"00787c04",
  2298 => x"447c3800",
  2299 => x"00387c44",
  2300 => x"24fcfc00",
  2301 => x"00183c24",
  2302 => x"243c1800",
  2303 => x"00fcfc24",
  2304 => x"047c7c00",
  2305 => x"00080c04",
  2306 => x"545c4800",
  2307 => x"00207454",
  2308 => x"7f3f0400",
  2309 => x"00004444",
  2310 => x"407c3c00",
  2311 => x"007c7c40",
  2312 => x"603c1c00",
  2313 => x"001c3c60",
  2314 => x"30607c3c",
  2315 => x"003c7c60",
  2316 => x"10386c44",
  2317 => x"00446c38",
  2318 => x"e0bc1c00",
  2319 => x"001c3c60",
  2320 => x"74644400",
  2321 => x"00444c5c",
  2322 => x"3e080800",
  2323 => x"00414177",
  2324 => x"7f000000",
  2325 => x"0000007f",
  2326 => x"77414100",
  2327 => x"0008083e",
  2328 => x"03010102",
  2329 => x"00010202",
  2330 => x"7f7f7f7f",
  2331 => x"007f7f7f",
  2332 => x"1c1c0808",
  2333 => x"7f7f3e3e",
  2334 => x"3e3e7f7f",
  2335 => x"08081c1c",
  2336 => x"7c181000",
  2337 => x"0010187c",
  2338 => x"7c301000",
  2339 => x"0010307c",
  2340 => x"60603010",
  2341 => x"00061e78",
  2342 => x"183c6642",
  2343 => x"0042663c",
  2344 => x"c26a3878",
  2345 => x"00386cc6",
  2346 => x"60000060",
  2347 => x"00600000",
  2348 => x"5c5b5e0e",
  2349 => x"86fc0e5d",
  2350 => x"fcc27e71",
  2351 => x"c04cbfe8",
  2352 => x"c41ec04b",
  2353 => x"c402ab66",
  2354 => x"c24dc087",
  2355 => x"754dc187",
  2356 => x"ee49731e",
  2357 => x"86c887e3",
  2358 => x"ef49e0c0",
  2359 => x"a4c487ec",
  2360 => x"f0496a4a",
  2361 => x"caf187f3",
  2362 => x"c184cc87",
  2363 => x"abb7c883",
  2364 => x"87cdff04",
  2365 => x"4d268efc",
  2366 => x"4b264c26",
  2367 => x"711e4f26",
  2368 => x"ecfcc24a",
  2369 => x"ecfcc25a",
  2370 => x"4978c748",
  2371 => x"2687e1fe",
  2372 => x"1e731e4f",
  2373 => x"b7c04a71",
  2374 => x"87d303aa",
  2375 => x"bff4e0c2",
  2376 => x"c187c405",
  2377 => x"c087c24b",
  2378 => x"f8e0c24b",
  2379 => x"c287c45b",
  2380 => x"fc5af8e0",
  2381 => x"f4e0c248",
  2382 => x"c14a78bf",
  2383 => x"a2c0c19a",
  2384 => x"87e8ec49",
  2385 => x"4f264b26",
  2386 => x"c44a711e",
  2387 => x"49721e66",
  2388 => x"fc87e0eb",
  2389 => x"1e4f268e",
  2390 => x"c348d4ff",
  2391 => x"d0ff78ff",
  2392 => x"78e1c048",
  2393 => x"c148d4ff",
  2394 => x"c4487178",
  2395 => x"08d4ff30",
  2396 => x"48d0ff78",
  2397 => x"2678e0c0",
  2398 => x"5b5e0e4f",
  2399 => x"f00e5d5c",
  2400 => x"48a6c886",
  2401 => x"ec4d78c0",
  2402 => x"80fc7ebf",
  2403 => x"bfe8fcc2",
  2404 => x"4cbfe878",
  2405 => x"bff4e0c2",
  2406 => x"87dde349",
  2407 => x"ca49eecb",
  2408 => x"4b7087d6",
  2409 => x"d2e749c7",
  2410 => x"05987087",
  2411 => x"496e87c8",
  2412 => x"c10299c1",
  2413 => x"4dc187c1",
  2414 => x"c27ebfec",
  2415 => x"49bff4e0",
  2416 => x"7387f6e2",
  2417 => x"87fcc949",
  2418 => x"d7029870",
  2419 => x"ece0c287",
  2420 => x"b9c149bf",
  2421 => x"59f0e0c2",
  2422 => x"87fbfd71",
  2423 => x"c949eecb",
  2424 => x"4b7087d6",
  2425 => x"d2e649c7",
  2426 => x"05987087",
  2427 => x"6e87c7ff",
  2428 => x"0599c149",
  2429 => x"7587fffe",
  2430 => x"e3c0029d",
  2431 => x"f4e0c287",
  2432 => x"bac14abf",
  2433 => x"5af8e0c2",
  2434 => x"0a7a0afc",
  2435 => x"c0c19ac1",
  2436 => x"d7e949a2",
  2437 => x"49dac187",
  2438 => x"c887e0e5",
  2439 => x"78c148a6",
  2440 => x"bff4e0c2",
  2441 => x"87e9c005",
  2442 => x"ffc34974",
  2443 => x"c01e7199",
  2444 => x"87d4fc49",
  2445 => x"b7c84974",
  2446 => x"c11e7129",
  2447 => x"87c8fc49",
  2448 => x"fdc386c8",
  2449 => x"87f3e449",
  2450 => x"e449fac3",
  2451 => x"d1c787ed",
  2452 => x"c3497487",
  2453 => x"b7c899ff",
  2454 => x"74b4712c",
  2455 => x"87df029c",
  2456 => x"bff0e0c2",
  2457 => x"87dcc749",
  2458 => x"c0059870",
  2459 => x"4cc087c4",
  2460 => x"e0c287d3",
  2461 => x"87c0c749",
  2462 => x"58f4e0c2",
  2463 => x"c287c6c0",
  2464 => x"c048f0e0",
  2465 => x"c8497478",
  2466 => x"87ce0599",
  2467 => x"e349f5c3",
  2468 => x"497087e9",
  2469 => x"c00299c2",
  2470 => x"fcc287e9",
  2471 => x"c002bfec",
  2472 => x"c14887c9",
  2473 => x"f0fcc288",
  2474 => x"c487d358",
  2475 => x"e0c14866",
  2476 => x"6e7e7080",
  2477 => x"c5c002bf",
  2478 => x"49ff4b87",
  2479 => x"a6c80f73",
  2480 => x"7478c148",
  2481 => x"0599c449",
  2482 => x"c387cec0",
  2483 => x"eae249f2",
  2484 => x"c2497087",
  2485 => x"f0c00299",
  2486 => x"ecfcc287",
  2487 => x"c7487ebf",
  2488 => x"c003a8b7",
  2489 => x"486e87cb",
  2490 => x"fcc280c1",
  2491 => x"d3c058f0",
  2492 => x"4866c487",
  2493 => x"7080e0c1",
  2494 => x"02bf6e7e",
  2495 => x"4b87c5c0",
  2496 => x"0f7349fe",
  2497 => x"c148a6c8",
  2498 => x"49fdc378",
  2499 => x"7087ece1",
  2500 => x"0299c249",
  2501 => x"c287e9c0",
  2502 => x"02bfecfc",
  2503 => x"c287c9c0",
  2504 => x"c048ecfc",
  2505 => x"87d3c078",
  2506 => x"c14866c4",
  2507 => x"7e7080e0",
  2508 => x"c002bf6e",
  2509 => x"fd4b87c5",
  2510 => x"c80f7349",
  2511 => x"78c148a6",
  2512 => x"e049fac3",
  2513 => x"497087f5",
  2514 => x"c00299c2",
  2515 => x"fcc287ea",
  2516 => x"c748bfec",
  2517 => x"c003a8b7",
  2518 => x"fcc287c9",
  2519 => x"78c748ec",
  2520 => x"c487d0c0",
  2521 => x"e0c14a66",
  2522 => x"c0026a82",
  2523 => x"fc4b87c5",
  2524 => x"c80f7349",
  2525 => x"78c148a6",
  2526 => x"fcc24dc0",
  2527 => x"50c048e4",
  2528 => x"c249eecb",
  2529 => x"4b7087f2",
  2530 => x"97e4fcc2",
  2531 => x"ddc105bf",
  2532 => x"c3497487",
  2533 => x"c00599f0",
  2534 => x"dac187cd",
  2535 => x"dadfff49",
  2536 => x"02987087",
  2537 => x"c187c7c1",
  2538 => x"4cbfe84d",
  2539 => x"99ffc349",
  2540 => x"712cb7c8",
  2541 => x"f4e0c2b4",
  2542 => x"daff49bf",
  2543 => x"497387fb",
  2544 => x"7087c1c2",
  2545 => x"c6c00298",
  2546 => x"e4fcc287",
  2547 => x"c250c148",
  2548 => x"bf97e4fc",
  2549 => x"87d6c005",
  2550 => x"f0c34974",
  2551 => x"c6ff0599",
  2552 => x"49dac187",
  2553 => x"87d3deff",
  2554 => x"fe059870",
  2555 => x"9d7587f9",
  2556 => x"87e0c002",
  2557 => x"c248a6cc",
  2558 => x"78bfecfc",
  2559 => x"cc4966cc",
  2560 => x"4866c491",
  2561 => x"7e708071",
  2562 => x"c002bf6e",
  2563 => x"cc4b87c6",
  2564 => x"0f734966",
  2565 => x"c00266c8",
  2566 => x"fcc287c8",
  2567 => x"f249bfec",
  2568 => x"8ef087ce",
  2569 => x"4c264d26",
  2570 => x"4f264b26",
  2571 => x"00000000",
  2572 => x"00000000",
  2573 => x"00000000",
  2574 => x"ff4a711e",
  2575 => x"7249bfc8",
  2576 => x"4f2648a1",
  2577 => x"bfc8ff1e",
  2578 => x"c0c0fe89",
  2579 => x"a9c0c0c0",
  2580 => x"c087c401",
  2581 => x"c187c24a",
  2582 => x"2648724a",
  2583 => x"5b5e0e4f",
  2584 => x"710e5d5c",
  2585 => x"4cd4ff4b",
  2586 => x"c04866d0",
  2587 => x"ff49d678",
  2588 => x"c387c5de",
  2589 => x"496c7cff",
  2590 => x"7199ffc3",
  2591 => x"f0c3494d",
  2592 => x"a9e0c199",
  2593 => x"c387cb05",
  2594 => x"486c7cff",
  2595 => x"66d098c3",
  2596 => x"ffc37808",
  2597 => x"494a6c7c",
  2598 => x"ffc331c8",
  2599 => x"714a6c7c",
  2600 => x"c84972b2",
  2601 => x"7cffc331",
  2602 => x"b2714a6c",
  2603 => x"31c84972",
  2604 => x"6c7cffc3",
  2605 => x"ffb2714a",
  2606 => x"e0c048d0",
  2607 => x"029b7378",
  2608 => x"7b7287c2",
  2609 => x"4d264875",
  2610 => x"4b264c26",
  2611 => x"261e4f26",
  2612 => x"5b5e0e4f",
  2613 => x"86f80e5c",
  2614 => x"a6c81e76",
  2615 => x"87fdfd49",
  2616 => x"4b7086c4",
  2617 => x"a8c4486e",
  2618 => x"87f4c203",
  2619 => x"f0c34a73",
  2620 => x"aad0c19a",
  2621 => x"c187c702",
  2622 => x"c205aae0",
  2623 => x"497387e2",
  2624 => x"c30299c8",
  2625 => x"87c6ff87",
  2626 => x"9cc34c73",
  2627 => x"c105acc2",
  2628 => x"66c487c4",
  2629 => x"7131c949",
  2630 => x"4a66c41e",
  2631 => x"c292c8c1",
  2632 => x"7249f0fc",
  2633 => x"c3ccfe81",
  2634 => x"ff49d887",
  2635 => x"c887c9db",
  2636 => x"eac21ec0",
  2637 => x"e2fd49d4",
  2638 => x"d0ff87c2",
  2639 => x"78e0c048",
  2640 => x"1ed4eac2",
  2641 => x"c14a66cc",
  2642 => x"fcc292c8",
  2643 => x"817249f0",
  2644 => x"87d2c7fe",
  2645 => x"acc186cc",
  2646 => x"87c4c105",
  2647 => x"c94966c4",
  2648 => x"c41e7131",
  2649 => x"c8c14a66",
  2650 => x"f0fcc292",
  2651 => x"fe817249",
  2652 => x"c287f9ca",
  2653 => x"c81ed4ea",
  2654 => x"c8c14a66",
  2655 => x"f0fcc292",
  2656 => x"fe817249",
  2657 => x"d787d0c5",
  2658 => x"ebd9ff49",
  2659 => x"1ec0c887",
  2660 => x"49d4eac2",
  2661 => x"87c1e0fd",
  2662 => x"d0ff86cc",
  2663 => x"78e0c048",
  2664 => x"4c268ef8",
  2665 => x"4f264b26",
  2666 => x"5c5b5e0e",
  2667 => x"86fc0e5d",
  2668 => x"d4ff4d71",
  2669 => x"7e66d44c",
  2670 => x"a8b7c348",
  2671 => x"87e3c101",
  2672 => x"66c41e75",
  2673 => x"93c8c14b",
  2674 => x"83f0fcc2",
  2675 => x"fefd4973",
  2676 => x"a3c887c7",
  2677 => x"ff496949",
  2678 => x"e1c848d0",
  2679 => x"717cdd78",
  2680 => x"98ffc348",
  2681 => x"4a717c70",
  2682 => x"722ab7c8",
  2683 => x"98ffc348",
  2684 => x"4a717c70",
  2685 => x"722ab7d0",
  2686 => x"98ffc348",
  2687 => x"48717c70",
  2688 => x"7028b7d8",
  2689 => x"7c7cc07c",
  2690 => x"7c7c7c7c",
  2691 => x"7c7c7c7c",
  2692 => x"d0ff7c7c",
  2693 => x"78e0c048",
  2694 => x"dc1e66c4",
  2695 => x"fcd7ff49",
  2696 => x"fc86c887",
  2697 => x"264d268e",
  2698 => x"264b264c",
  2699 => x"1ec01e4f",
  2700 => x"bfc8e9c2",
  2701 => x"87f0fd49",
  2702 => x"bfcce9c2",
  2703 => x"e5dcfe49",
  2704 => x"fc48c087",
  2705 => x"004f268e",
  2706 => x"00002a50",
  2707 => x"00002a5c",
  2708 => x"3834585a",
  2709 => x"20202020",
  2710 => x"00444856",
  2711 => x"3834585a",
  2712 => x"20202020",
  2713 => x"004d4f52",
  2714 => x"00001d8f",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
