
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom2 is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom2 is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"08",x"d4",x"ff",x"48"),
     1 => (x"1e",x"4f",x"26",x"78"),
     2 => (x"c8",x"48",x"d0",x"ff"),
     3 => (x"48",x"71",x"78",x"e1"),
     4 => (x"78",x"08",x"d4",x"ff"),
     5 => (x"ff",x"48",x"66",x"c4"),
     6 => (x"26",x"78",x"08",x"d4"),
     7 => (x"4a",x"71",x"1e",x"4f"),
     8 => (x"1e",x"49",x"66",x"c4"),
     9 => (x"de",x"ff",x"49",x"72"),
    10 => (x"48",x"d0",x"ff",x"87"),
    11 => (x"fc",x"78",x"e0",x"c0"),
    12 => (x"1e",x"4f",x"26",x"8e"),
    13 => (x"4a",x"71",x"1e",x"73"),
    14 => (x"ab",x"b7",x"c2",x"4b"),
    15 => (x"a3",x"87",x"c8",x"03"),
    16 => (x"ff",x"c3",x"4a",x"49"),
    17 => (x"ce",x"87",x"c7",x"9a"),
    18 => (x"c3",x"4a",x"49",x"a3"),
    19 => (x"66",x"c8",x"9a",x"ff"),
    20 => (x"49",x"72",x"1e",x"49"),
    21 => (x"fc",x"87",x"c6",x"ff"),
    22 => (x"26",x"4b",x"26",x"8e"),
    23 => (x"d0",x"ff",x"1e",x"4f"),
    24 => (x"78",x"c9",x"c8",x"48"),
    25 => (x"d4",x"ff",x"48",x"71"),
    26 => (x"4f",x"26",x"78",x"08"),
    27 => (x"49",x"4a",x"71",x"1e"),
    28 => (x"d0",x"ff",x"87",x"eb"),
    29 => (x"26",x"78",x"c8",x"48"),
    30 => (x"1e",x"73",x"1e",x"4f"),
    31 => (x"fc",x"c2",x"4b",x"71"),
    32 => (x"c3",x"02",x"bf",x"e0"),
    33 => (x"87",x"eb",x"c2",x"87"),
    34 => (x"c8",x"48",x"d0",x"ff"),
    35 => (x"48",x"73",x"78",x"c9"),
    36 => (x"ff",x"b0",x"e0",x"c0"),
    37 => (x"c2",x"78",x"08",x"d4"),
    38 => (x"c0",x"48",x"d4",x"fc"),
    39 => (x"02",x"66",x"c8",x"78"),
    40 => (x"ff",x"c3",x"87",x"c5"),
    41 => (x"c0",x"87",x"c2",x"49"),
    42 => (x"dc",x"fc",x"c2",x"49"),
    43 => (x"02",x"66",x"cc",x"59"),
    44 => (x"d5",x"c5",x"87",x"c6"),
    45 => (x"87",x"c4",x"4a",x"d5"),
    46 => (x"4a",x"ff",x"ff",x"cf"),
    47 => (x"5a",x"e0",x"fc",x"c2"),
    48 => (x"48",x"e0",x"fc",x"c2"),
    49 => (x"4b",x"26",x"78",x"c1"),
    50 => (x"5e",x"0e",x"4f",x"26"),
    51 => (x"0e",x"5d",x"5c",x"5b"),
    52 => (x"fc",x"c2",x"4d",x"71"),
    53 => (x"75",x"4b",x"bf",x"dc"),
    54 => (x"87",x"cb",x"02",x"9d"),
    55 => (x"c2",x"91",x"c8",x"49"),
    56 => (x"71",x"4a",x"f0",x"c1"),
    57 => (x"c2",x"87",x"c4",x"82"),
    58 => (x"c0",x"4a",x"f0",x"c5"),
    59 => (x"73",x"49",x"12",x"4c"),
    60 => (x"d8",x"fc",x"c2",x"99"),
    61 => (x"b8",x"71",x"48",x"bf"),
    62 => (x"78",x"08",x"d4",x"ff"),
    63 => (x"84",x"2b",x"b7",x"c1"),
    64 => (x"04",x"ac",x"b7",x"c8"),
    65 => (x"fc",x"c2",x"87",x"e7"),
    66 => (x"c8",x"48",x"bf",x"d4"),
    67 => (x"d8",x"fc",x"c2",x"80"),
    68 => (x"26",x"4d",x"26",x"58"),
    69 => (x"26",x"4b",x"26",x"4c"),
    70 => (x"1e",x"73",x"1e",x"4f"),
    71 => (x"4a",x"13",x"4b",x"71"),
    72 => (x"87",x"cb",x"02",x"9a"),
    73 => (x"e1",x"fe",x"49",x"72"),
    74 => (x"9a",x"4a",x"13",x"87"),
    75 => (x"26",x"87",x"f5",x"05"),
    76 => (x"1e",x"4f",x"26",x"4b"),
    77 => (x"bf",x"d4",x"fc",x"c2"),
    78 => (x"d4",x"fc",x"c2",x"49"),
    79 => (x"78",x"a1",x"c1",x"48"),
    80 => (x"a9",x"b7",x"c0",x"c4"),
    81 => (x"ff",x"87",x"db",x"03"),
    82 => (x"fc",x"c2",x"48",x"d4"),
    83 => (x"c2",x"78",x"bf",x"d8"),
    84 => (x"49",x"bf",x"d4",x"fc"),
    85 => (x"48",x"d4",x"fc",x"c2"),
    86 => (x"c4",x"78",x"a1",x"c1"),
    87 => (x"04",x"a9",x"b7",x"c0"),
    88 => (x"d0",x"ff",x"87",x"e5"),
    89 => (x"c2",x"78",x"c8",x"48"),
    90 => (x"c0",x"48",x"e0",x"fc"),
    91 => (x"00",x"4f",x"26",x"78"),
    92 => (x"00",x"00",x"00",x"00"),
    93 => (x"00",x"00",x"00",x"00"),
    94 => (x"5f",x"00",x"00",x"00"),
    95 => (x"00",x"00",x"00",x"5f"),
    96 => (x"00",x"03",x"03",x"00"),
    97 => (x"00",x"00",x"03",x"03"),
    98 => (x"14",x"7f",x"7f",x"14"),
    99 => (x"00",x"14",x"7f",x"7f"),
   100 => (x"6b",x"2e",x"24",x"00"),
   101 => (x"00",x"12",x"3a",x"6b"),
   102 => (x"18",x"36",x"6a",x"4c"),
   103 => (x"00",x"32",x"56",x"6c"),
   104 => (x"59",x"4f",x"7e",x"30"),
   105 => (x"40",x"68",x"3a",x"77"),
   106 => (x"07",x"04",x"00",x"00"),
   107 => (x"00",x"00",x"00",x"03"),
   108 => (x"3e",x"1c",x"00",x"00"),
   109 => (x"00",x"00",x"41",x"63"),
   110 => (x"63",x"41",x"00",x"00"),
   111 => (x"00",x"00",x"1c",x"3e"),
   112 => (x"1c",x"3e",x"2a",x"08"),
   113 => (x"08",x"2a",x"3e",x"1c"),
   114 => (x"3e",x"08",x"08",x"00"),
   115 => (x"00",x"08",x"08",x"3e"),
   116 => (x"e0",x"80",x"00",x"00"),
   117 => (x"00",x"00",x"00",x"60"),
   118 => (x"08",x"08",x"08",x"00"),
   119 => (x"00",x"08",x"08",x"08"),
   120 => (x"60",x"00",x"00",x"00"),
   121 => (x"00",x"00",x"00",x"60"),
   122 => (x"18",x"30",x"60",x"40"),
   123 => (x"01",x"03",x"06",x"0c"),
   124 => (x"59",x"7f",x"3e",x"00"),
   125 => (x"00",x"3e",x"7f",x"4d"),
   126 => (x"7f",x"06",x"04",x"00"),
   127 => (x"00",x"00",x"00",x"7f"),
   128 => (x"71",x"63",x"42",x"00"),
   129 => (x"00",x"46",x"4f",x"59"),
   130 => (x"49",x"63",x"22",x"00"),
   131 => (x"00",x"36",x"7f",x"49"),
   132 => (x"13",x"16",x"1c",x"18"),
   133 => (x"00",x"10",x"7f",x"7f"),
   134 => (x"45",x"67",x"27",x"00"),
   135 => (x"00",x"39",x"7d",x"45"),
   136 => (x"4b",x"7e",x"3c",x"00"),
   137 => (x"00",x"30",x"79",x"49"),
   138 => (x"71",x"01",x"01",x"00"),
   139 => (x"00",x"07",x"0f",x"79"),
   140 => (x"49",x"7f",x"36",x"00"),
   141 => (x"00",x"36",x"7f",x"49"),
   142 => (x"49",x"4f",x"06",x"00"),
   143 => (x"00",x"1e",x"3f",x"69"),
   144 => (x"66",x"00",x"00",x"00"),
   145 => (x"00",x"00",x"00",x"66"),
   146 => (x"e6",x"80",x"00",x"00"),
   147 => (x"00",x"00",x"00",x"66"),
   148 => (x"14",x"08",x"08",x"00"),
   149 => (x"00",x"22",x"22",x"14"),
   150 => (x"14",x"14",x"14",x"00"),
   151 => (x"00",x"14",x"14",x"14"),
   152 => (x"14",x"22",x"22",x"00"),
   153 => (x"00",x"08",x"08",x"14"),
   154 => (x"51",x"03",x"02",x"00"),
   155 => (x"00",x"06",x"0f",x"59"),
   156 => (x"5d",x"41",x"7f",x"3e"),
   157 => (x"00",x"1e",x"1f",x"55"),
   158 => (x"09",x"7f",x"7e",x"00"),
   159 => (x"00",x"7e",x"7f",x"09"),
   160 => (x"49",x"7f",x"7f",x"00"),
   161 => (x"00",x"36",x"7f",x"49"),
   162 => (x"63",x"3e",x"1c",x"00"),
   163 => (x"00",x"41",x"41",x"41"),
   164 => (x"41",x"7f",x"7f",x"00"),
   165 => (x"00",x"1c",x"3e",x"63"),
   166 => (x"49",x"7f",x"7f",x"00"),
   167 => (x"00",x"41",x"41",x"49"),
   168 => (x"09",x"7f",x"7f",x"00"),
   169 => (x"00",x"01",x"01",x"09"),
   170 => (x"41",x"7f",x"3e",x"00"),
   171 => (x"00",x"7a",x"7b",x"49"),
   172 => (x"08",x"7f",x"7f",x"00"),
   173 => (x"00",x"7f",x"7f",x"08"),
   174 => (x"7f",x"41",x"00",x"00"),
   175 => (x"00",x"00",x"41",x"7f"),
   176 => (x"40",x"60",x"20",x"00"),
   177 => (x"00",x"3f",x"7f",x"40"),
   178 => (x"1c",x"08",x"7f",x"7f"),
   179 => (x"00",x"41",x"63",x"36"),
   180 => (x"40",x"7f",x"7f",x"00"),
   181 => (x"00",x"40",x"40",x"40"),
   182 => (x"0c",x"06",x"7f",x"7f"),
   183 => (x"00",x"7f",x"7f",x"06"),
   184 => (x"0c",x"06",x"7f",x"7f"),
   185 => (x"00",x"7f",x"7f",x"18"),
   186 => (x"41",x"7f",x"3e",x"00"),
   187 => (x"00",x"3e",x"7f",x"41"),
   188 => (x"09",x"7f",x"7f",x"00"),
   189 => (x"00",x"06",x"0f",x"09"),
   190 => (x"61",x"41",x"7f",x"3e"),
   191 => (x"00",x"40",x"7e",x"7f"),
   192 => (x"09",x"7f",x"7f",x"00"),
   193 => (x"00",x"66",x"7f",x"19"),
   194 => (x"4d",x"6f",x"26",x"00"),
   195 => (x"00",x"32",x"7b",x"59"),
   196 => (x"7f",x"01",x"01",x"00"),
   197 => (x"00",x"01",x"01",x"7f"),
   198 => (x"40",x"7f",x"3f",x"00"),
   199 => (x"00",x"3f",x"7f",x"40"),
   200 => (x"70",x"3f",x"0f",x"00"),
   201 => (x"00",x"0f",x"3f",x"70"),
   202 => (x"18",x"30",x"7f",x"7f"),
   203 => (x"00",x"7f",x"7f",x"30"),
   204 => (x"1c",x"36",x"63",x"41"),
   205 => (x"41",x"63",x"36",x"1c"),
   206 => (x"7c",x"06",x"03",x"01"),
   207 => (x"01",x"03",x"06",x"7c"),
   208 => (x"4d",x"59",x"71",x"61"),
   209 => (x"00",x"41",x"43",x"47"),
   210 => (x"7f",x"7f",x"00",x"00"),
   211 => (x"00",x"00",x"41",x"41"),
   212 => (x"0c",x"06",x"03",x"01"),
   213 => (x"40",x"60",x"30",x"18"),
   214 => (x"41",x"41",x"00",x"00"),
   215 => (x"00",x"00",x"7f",x"7f"),
   216 => (x"03",x"06",x"0c",x"08"),
   217 => (x"00",x"08",x"0c",x"06"),
   218 => (x"80",x"80",x"80",x"80"),
   219 => (x"00",x"80",x"80",x"80"),
   220 => (x"03",x"00",x"00",x"00"),
   221 => (x"00",x"00",x"04",x"07"),
   222 => (x"54",x"74",x"20",x"00"),
   223 => (x"00",x"78",x"7c",x"54"),
   224 => (x"44",x"7f",x"7f",x"00"),
   225 => (x"00",x"38",x"7c",x"44"),
   226 => (x"44",x"7c",x"38",x"00"),
   227 => (x"00",x"00",x"44",x"44"),
   228 => (x"44",x"7c",x"38",x"00"),
   229 => (x"00",x"7f",x"7f",x"44"),
   230 => (x"54",x"7c",x"38",x"00"),
   231 => (x"00",x"18",x"5c",x"54"),
   232 => (x"7f",x"7e",x"04",x"00"),
   233 => (x"00",x"00",x"05",x"05"),
   234 => (x"a4",x"bc",x"18",x"00"),
   235 => (x"00",x"7c",x"fc",x"a4"),
   236 => (x"04",x"7f",x"7f",x"00"),
   237 => (x"00",x"78",x"7c",x"04"),
   238 => (x"3d",x"00",x"00",x"00"),
   239 => (x"00",x"00",x"40",x"7d"),
   240 => (x"80",x"80",x"80",x"00"),
   241 => (x"00",x"00",x"7d",x"fd"),
   242 => (x"10",x"7f",x"7f",x"00"),
   243 => (x"00",x"44",x"6c",x"38"),
   244 => (x"3f",x"00",x"00",x"00"),
   245 => (x"00",x"00",x"40",x"7f"),
   246 => (x"18",x"0c",x"7c",x"7c"),
   247 => (x"00",x"78",x"7c",x"0c"),
   248 => (x"04",x"7c",x"7c",x"00"),
   249 => (x"00",x"78",x"7c",x"04"),
   250 => (x"44",x"7c",x"38",x"00"),
   251 => (x"00",x"38",x"7c",x"44"),
   252 => (x"24",x"fc",x"fc",x"00"),
   253 => (x"00",x"18",x"3c",x"24"),
   254 => (x"24",x"3c",x"18",x"00"),
   255 => (x"00",x"fc",x"fc",x"24"),
   256 => (x"04",x"7c",x"7c",x"00"),
   257 => (x"00",x"08",x"0c",x"04"),
   258 => (x"54",x"5c",x"48",x"00"),
   259 => (x"00",x"20",x"74",x"54"),
   260 => (x"7f",x"3f",x"04",x"00"),
   261 => (x"00",x"00",x"44",x"44"),
   262 => (x"40",x"7c",x"3c",x"00"),
   263 => (x"00",x"7c",x"7c",x"40"),
   264 => (x"60",x"3c",x"1c",x"00"),
   265 => (x"00",x"1c",x"3c",x"60"),
   266 => (x"30",x"60",x"7c",x"3c"),
   267 => (x"00",x"3c",x"7c",x"60"),
   268 => (x"10",x"38",x"6c",x"44"),
   269 => (x"00",x"44",x"6c",x"38"),
   270 => (x"e0",x"bc",x"1c",x"00"),
   271 => (x"00",x"1c",x"3c",x"60"),
   272 => (x"74",x"64",x"44",x"00"),
   273 => (x"00",x"44",x"4c",x"5c"),
   274 => (x"3e",x"08",x"08",x"00"),
   275 => (x"00",x"41",x"41",x"77"),
   276 => (x"7f",x"00",x"00",x"00"),
   277 => (x"00",x"00",x"00",x"7f"),
   278 => (x"77",x"41",x"41",x"00"),
   279 => (x"00",x"08",x"08",x"3e"),
   280 => (x"03",x"01",x"01",x"02"),
   281 => (x"00",x"01",x"02",x"02"),
   282 => (x"7f",x"7f",x"7f",x"7f"),
   283 => (x"00",x"7f",x"7f",x"7f"),
   284 => (x"1c",x"1c",x"08",x"08"),
   285 => (x"7f",x"7f",x"3e",x"3e"),
   286 => (x"3e",x"3e",x"7f",x"7f"),
   287 => (x"08",x"08",x"1c",x"1c"),
   288 => (x"7c",x"18",x"10",x"00"),
   289 => (x"00",x"10",x"18",x"7c"),
   290 => (x"7c",x"30",x"10",x"00"),
   291 => (x"00",x"10",x"30",x"7c"),
   292 => (x"60",x"60",x"30",x"10"),
   293 => (x"00",x"06",x"1e",x"78"),
   294 => (x"18",x"3c",x"66",x"42"),
   295 => (x"00",x"42",x"66",x"3c"),
   296 => (x"c2",x"6a",x"38",x"78"),
   297 => (x"00",x"38",x"6c",x"c6"),
   298 => (x"60",x"00",x"00",x"60"),
   299 => (x"00",x"60",x"00",x"00"),
   300 => (x"5c",x"5b",x"5e",x"0e"),
   301 => (x"86",x"fc",x"0e",x"5d"),
   302 => (x"fc",x"c2",x"7e",x"71"),
   303 => (x"c0",x"4c",x"bf",x"e8"),
   304 => (x"c4",x"1e",x"c0",x"4b"),
   305 => (x"c4",x"02",x"ab",x"66"),
   306 => (x"c2",x"4d",x"c0",x"87"),
   307 => (x"75",x"4d",x"c1",x"87"),
   308 => (x"ee",x"49",x"73",x"1e"),
   309 => (x"86",x"c8",x"87",x"e3"),
   310 => (x"ef",x"49",x"e0",x"c0"),
   311 => (x"a4",x"c4",x"87",x"ec"),
   312 => (x"f0",x"49",x"6a",x"4a"),
   313 => (x"ca",x"f1",x"87",x"f3"),
   314 => (x"c1",x"84",x"cc",x"87"),
   315 => (x"ab",x"b7",x"c8",x"83"),
   316 => (x"87",x"cd",x"ff",x"04"),
   317 => (x"4d",x"26",x"8e",x"fc"),
   318 => (x"4b",x"26",x"4c",x"26"),
   319 => (x"71",x"1e",x"4f",x"26"),
   320 => (x"ec",x"fc",x"c2",x"4a"),
   321 => (x"ec",x"fc",x"c2",x"5a"),
   322 => (x"49",x"78",x"c7",x"48"),
   323 => (x"26",x"87",x"e1",x"fe"),
   324 => (x"1e",x"73",x"1e",x"4f"),
   325 => (x"b7",x"c0",x"4a",x"71"),
   326 => (x"87",x"d3",x"03",x"aa"),
   327 => (x"bf",x"f4",x"e0",x"c2"),
   328 => (x"c1",x"87",x"c4",x"05"),
   329 => (x"c0",x"87",x"c2",x"4b"),
   330 => (x"f8",x"e0",x"c2",x"4b"),
   331 => (x"c2",x"87",x"c4",x"5b"),
   332 => (x"fc",x"5a",x"f8",x"e0"),
   333 => (x"f4",x"e0",x"c2",x"48"),
   334 => (x"c1",x"4a",x"78",x"bf"),
   335 => (x"a2",x"c0",x"c1",x"9a"),
   336 => (x"87",x"e8",x"ec",x"49"),
   337 => (x"4f",x"26",x"4b",x"26"),
   338 => (x"c4",x"4a",x"71",x"1e"),
   339 => (x"49",x"72",x"1e",x"66"),
   340 => (x"fc",x"87",x"e0",x"eb"),
   341 => (x"1e",x"4f",x"26",x"8e"),
   342 => (x"c3",x"48",x"d4",x"ff"),
   343 => (x"d0",x"ff",x"78",x"ff"),
   344 => (x"78",x"e1",x"c0",x"48"),
   345 => (x"c1",x"48",x"d4",x"ff"),
   346 => (x"c4",x"48",x"71",x"78"),
   347 => (x"08",x"d4",x"ff",x"30"),
   348 => (x"48",x"d0",x"ff",x"78"),
   349 => (x"26",x"78",x"e0",x"c0"),
   350 => (x"5b",x"5e",x"0e",x"4f"),
   351 => (x"f0",x"0e",x"5d",x"5c"),
   352 => (x"48",x"a6",x"c8",x"86"),
   353 => (x"ec",x"4d",x"78",x"c0"),
   354 => (x"80",x"fc",x"7e",x"bf"),
   355 => (x"bf",x"e8",x"fc",x"c2"),
   356 => (x"4c",x"bf",x"e8",x"78"),
   357 => (x"bf",x"f4",x"e0",x"c2"),
   358 => (x"87",x"dd",x"e3",x"49"),
   359 => (x"ca",x"49",x"ee",x"cb"),
   360 => (x"4b",x"70",x"87",x"d6"),
   361 => (x"d2",x"e7",x"49",x"c7"),
   362 => (x"05",x"98",x"70",x"87"),
   363 => (x"49",x"6e",x"87",x"c8"),
   364 => (x"c1",x"02",x"99",x"c1"),
   365 => (x"4d",x"c1",x"87",x"c1"),
   366 => (x"c2",x"7e",x"bf",x"ec"),
   367 => (x"49",x"bf",x"f4",x"e0"),
   368 => (x"73",x"87",x"f6",x"e2"),
   369 => (x"87",x"fc",x"c9",x"49"),
   370 => (x"d7",x"02",x"98",x"70"),
   371 => (x"ec",x"e0",x"c2",x"87"),
   372 => (x"b9",x"c1",x"49",x"bf"),
   373 => (x"59",x"f0",x"e0",x"c2"),
   374 => (x"87",x"fb",x"fd",x"71"),
   375 => (x"c9",x"49",x"ee",x"cb"),
   376 => (x"4b",x"70",x"87",x"d6"),
   377 => (x"d2",x"e6",x"49",x"c7"),
   378 => (x"05",x"98",x"70",x"87"),
   379 => (x"6e",x"87",x"c7",x"ff"),
   380 => (x"05",x"99",x"c1",x"49"),
   381 => (x"75",x"87",x"ff",x"fe"),
   382 => (x"e3",x"c0",x"02",x"9d"),
   383 => (x"f4",x"e0",x"c2",x"87"),
   384 => (x"ba",x"c1",x"4a",x"bf"),
   385 => (x"5a",x"f8",x"e0",x"c2"),
   386 => (x"0a",x"7a",x"0a",x"fc"),
   387 => (x"c0",x"c1",x"9a",x"c1"),
   388 => (x"d7",x"e9",x"49",x"a2"),
   389 => (x"49",x"da",x"c1",x"87"),
   390 => (x"c8",x"87",x"e0",x"e5"),
   391 => (x"78",x"c1",x"48",x"a6"),
   392 => (x"bf",x"f4",x"e0",x"c2"),
   393 => (x"87",x"e9",x"c0",x"05"),
   394 => (x"ff",x"c3",x"49",x"74"),
   395 => (x"c0",x"1e",x"71",x"99"),
   396 => (x"87",x"d4",x"fc",x"49"),
   397 => (x"b7",x"c8",x"49",x"74"),
   398 => (x"c1",x"1e",x"71",x"29"),
   399 => (x"87",x"c8",x"fc",x"49"),
   400 => (x"fd",x"c3",x"86",x"c8"),
   401 => (x"87",x"f3",x"e4",x"49"),
   402 => (x"e4",x"49",x"fa",x"c3"),
   403 => (x"d1",x"c7",x"87",x"ed"),
   404 => (x"c3",x"49",x"74",x"87"),
   405 => (x"b7",x"c8",x"99",x"ff"),
   406 => (x"74",x"b4",x"71",x"2c"),
   407 => (x"87",x"df",x"02",x"9c"),
   408 => (x"bf",x"f0",x"e0",x"c2"),
   409 => (x"87",x"dc",x"c7",x"49"),
   410 => (x"c0",x"05",x"98",x"70"),
   411 => (x"4c",x"c0",x"87",x"c4"),
   412 => (x"e0",x"c2",x"87",x"d3"),
   413 => (x"87",x"c0",x"c7",x"49"),
   414 => (x"58",x"f4",x"e0",x"c2"),
   415 => (x"c2",x"87",x"c6",x"c0"),
   416 => (x"c0",x"48",x"f0",x"e0"),
   417 => (x"c8",x"49",x"74",x"78"),
   418 => (x"87",x"ce",x"05",x"99"),
   419 => (x"e3",x"49",x"f5",x"c3"),
   420 => (x"49",x"70",x"87",x"e9"),
   421 => (x"c0",x"02",x"99",x"c2"),
   422 => (x"fc",x"c2",x"87",x"e9"),
   423 => (x"c0",x"02",x"bf",x"ec"),
   424 => (x"c1",x"48",x"87",x"c9"),
   425 => (x"f0",x"fc",x"c2",x"88"),
   426 => (x"c4",x"87",x"d3",x"58"),
   427 => (x"e0",x"c1",x"48",x"66"),
   428 => (x"6e",x"7e",x"70",x"80"),
   429 => (x"c5",x"c0",x"02",x"bf"),
   430 => (x"49",x"ff",x"4b",x"87"),
   431 => (x"a6",x"c8",x"0f",x"73"),
   432 => (x"74",x"78",x"c1",x"48"),
   433 => (x"05",x"99",x"c4",x"49"),
   434 => (x"c3",x"87",x"ce",x"c0"),
   435 => (x"ea",x"e2",x"49",x"f2"),
   436 => (x"c2",x"49",x"70",x"87"),
   437 => (x"f0",x"c0",x"02",x"99"),
   438 => (x"ec",x"fc",x"c2",x"87"),
   439 => (x"c7",x"48",x"7e",x"bf"),
   440 => (x"c0",x"03",x"a8",x"b7"),
   441 => (x"48",x"6e",x"87",x"cb"),
   442 => (x"fc",x"c2",x"80",x"c1"),
   443 => (x"d3",x"c0",x"58",x"f0"),
   444 => (x"48",x"66",x"c4",x"87"),
   445 => (x"70",x"80",x"e0",x"c1"),
   446 => (x"02",x"bf",x"6e",x"7e"),
   447 => (x"4b",x"87",x"c5",x"c0"),
   448 => (x"0f",x"73",x"49",x"fe"),
   449 => (x"c1",x"48",x"a6",x"c8"),
   450 => (x"49",x"fd",x"c3",x"78"),
   451 => (x"70",x"87",x"ec",x"e1"),
   452 => (x"02",x"99",x"c2",x"49"),
   453 => (x"c2",x"87",x"e9",x"c0"),
   454 => (x"02",x"bf",x"ec",x"fc"),
   455 => (x"c2",x"87",x"c9",x"c0"),
   456 => (x"c0",x"48",x"ec",x"fc"),
   457 => (x"87",x"d3",x"c0",x"78"),
   458 => (x"c1",x"48",x"66",x"c4"),
   459 => (x"7e",x"70",x"80",x"e0"),
   460 => (x"c0",x"02",x"bf",x"6e"),
   461 => (x"fd",x"4b",x"87",x"c5"),
   462 => (x"c8",x"0f",x"73",x"49"),
   463 => (x"78",x"c1",x"48",x"a6"),
   464 => (x"e0",x"49",x"fa",x"c3"),
   465 => (x"49",x"70",x"87",x"f5"),
   466 => (x"c0",x"02",x"99",x"c2"),
   467 => (x"fc",x"c2",x"87",x"ea"),
   468 => (x"c7",x"48",x"bf",x"ec"),
   469 => (x"c0",x"03",x"a8",x"b7"),
   470 => (x"fc",x"c2",x"87",x"c9"),
   471 => (x"78",x"c7",x"48",x"ec"),
   472 => (x"c4",x"87",x"d0",x"c0"),
   473 => (x"e0",x"c1",x"4a",x"66"),
   474 => (x"c0",x"02",x"6a",x"82"),
   475 => (x"fc",x"4b",x"87",x"c5"),
   476 => (x"c8",x"0f",x"73",x"49"),
   477 => (x"78",x"c1",x"48",x"a6"),
   478 => (x"fc",x"c2",x"4d",x"c0"),
   479 => (x"50",x"c0",x"48",x"e4"),
   480 => (x"c2",x"49",x"ee",x"cb"),
   481 => (x"4b",x"70",x"87",x"f2"),
   482 => (x"97",x"e4",x"fc",x"c2"),
   483 => (x"dd",x"c1",x"05",x"bf"),
   484 => (x"c3",x"49",x"74",x"87"),
   485 => (x"c0",x"05",x"99",x"f0"),
   486 => (x"da",x"c1",x"87",x"cd"),
   487 => (x"da",x"df",x"ff",x"49"),
   488 => (x"02",x"98",x"70",x"87"),
   489 => (x"c1",x"87",x"c7",x"c1"),
   490 => (x"4c",x"bf",x"e8",x"4d"),
   491 => (x"99",x"ff",x"c3",x"49"),
   492 => (x"71",x"2c",x"b7",x"c8"),
   493 => (x"f4",x"e0",x"c2",x"b4"),
   494 => (x"da",x"ff",x"49",x"bf"),
   495 => (x"49",x"73",x"87",x"fb"),
   496 => (x"70",x"87",x"c1",x"c2"),
   497 => (x"c6",x"c0",x"02",x"98"),
   498 => (x"e4",x"fc",x"c2",x"87"),
   499 => (x"c2",x"50",x"c1",x"48"),
   500 => (x"bf",x"97",x"e4",x"fc"),
   501 => (x"87",x"d6",x"c0",x"05"),
   502 => (x"f0",x"c3",x"49",x"74"),
   503 => (x"c6",x"ff",x"05",x"99"),
   504 => (x"49",x"da",x"c1",x"87"),
   505 => (x"87",x"d3",x"de",x"ff"),
   506 => (x"fe",x"05",x"98",x"70"),
   507 => (x"9d",x"75",x"87",x"f9"),
   508 => (x"87",x"e0",x"c0",x"02"),
   509 => (x"c2",x"48",x"a6",x"cc"),
   510 => (x"78",x"bf",x"ec",x"fc"),
   511 => (x"cc",x"49",x"66",x"cc"),
   512 => (x"48",x"66",x"c4",x"91"),
   513 => (x"7e",x"70",x"80",x"71"),
   514 => (x"c0",x"02",x"bf",x"6e"),
   515 => (x"cc",x"4b",x"87",x"c6"),
   516 => (x"0f",x"73",x"49",x"66"),
   517 => (x"c0",x"02",x"66",x"c8"),
   518 => (x"fc",x"c2",x"87",x"c8"),
   519 => (x"f2",x"49",x"bf",x"ec"),
   520 => (x"8e",x"f0",x"87",x"ce"),
   521 => (x"4c",x"26",x"4d",x"26"),
   522 => (x"4f",x"26",x"4b",x"26"),
   523 => (x"00",x"00",x"00",x"00"),
   524 => (x"00",x"00",x"00",x"00"),
   525 => (x"00",x"00",x"00",x"00"),
   526 => (x"ff",x"4a",x"71",x"1e"),
   527 => (x"72",x"49",x"bf",x"c8"),
   528 => (x"4f",x"26",x"48",x"a1"),
   529 => (x"bf",x"c8",x"ff",x"1e"),
   530 => (x"c0",x"c0",x"fe",x"89"),
   531 => (x"a9",x"c0",x"c0",x"c0"),
   532 => (x"c0",x"87",x"c4",x"01"),
   533 => (x"c1",x"87",x"c2",x"4a"),
   534 => (x"26",x"48",x"72",x"4a"),
   535 => (x"5b",x"5e",x"0e",x"4f"),
   536 => (x"71",x"0e",x"5d",x"5c"),
   537 => (x"4c",x"d4",x"ff",x"4b"),
   538 => (x"c0",x"48",x"66",x"d0"),
   539 => (x"ff",x"49",x"d6",x"78"),
   540 => (x"c3",x"87",x"c5",x"de"),
   541 => (x"49",x"6c",x"7c",x"ff"),
   542 => (x"71",x"99",x"ff",x"c3"),
   543 => (x"f0",x"c3",x"49",x"4d"),
   544 => (x"a9",x"e0",x"c1",x"99"),
   545 => (x"c3",x"87",x"cb",x"05"),
   546 => (x"48",x"6c",x"7c",x"ff"),
   547 => (x"66",x"d0",x"98",x"c3"),
   548 => (x"ff",x"c3",x"78",x"08"),
   549 => (x"49",x"4a",x"6c",x"7c"),
   550 => (x"ff",x"c3",x"31",x"c8"),
   551 => (x"71",x"4a",x"6c",x"7c"),
   552 => (x"c8",x"49",x"72",x"b2"),
   553 => (x"7c",x"ff",x"c3",x"31"),
   554 => (x"b2",x"71",x"4a",x"6c"),
   555 => (x"31",x"c8",x"49",x"72"),
   556 => (x"6c",x"7c",x"ff",x"c3"),
   557 => (x"ff",x"b2",x"71",x"4a"),
   558 => (x"e0",x"c0",x"48",x"d0"),
   559 => (x"02",x"9b",x"73",x"78"),
   560 => (x"7b",x"72",x"87",x"c2"),
   561 => (x"4d",x"26",x"48",x"75"),
   562 => (x"4b",x"26",x"4c",x"26"),
   563 => (x"26",x"1e",x"4f",x"26"),
   564 => (x"5b",x"5e",x"0e",x"4f"),
   565 => (x"86",x"f8",x"0e",x"5c"),
   566 => (x"a6",x"c8",x"1e",x"76"),
   567 => (x"87",x"fd",x"fd",x"49"),
   568 => (x"4b",x"70",x"86",x"c4"),
   569 => (x"a8",x"c4",x"48",x"6e"),
   570 => (x"87",x"f4",x"c2",x"03"),
   571 => (x"f0",x"c3",x"4a",x"73"),
   572 => (x"aa",x"d0",x"c1",x"9a"),
   573 => (x"c1",x"87",x"c7",x"02"),
   574 => (x"c2",x"05",x"aa",x"e0"),
   575 => (x"49",x"73",x"87",x"e2"),
   576 => (x"c3",x"02",x"99",x"c8"),
   577 => (x"87",x"c6",x"ff",x"87"),
   578 => (x"9c",x"c3",x"4c",x"73"),
   579 => (x"c1",x"05",x"ac",x"c2"),
   580 => (x"66",x"c4",x"87",x"c4"),
   581 => (x"71",x"31",x"c9",x"49"),
   582 => (x"4a",x"66",x"c4",x"1e"),
   583 => (x"c2",x"92",x"c8",x"c1"),
   584 => (x"72",x"49",x"f0",x"fc"),
   585 => (x"c3",x"cc",x"fe",x"81"),
   586 => (x"ff",x"49",x"d8",x"87"),
   587 => (x"c8",x"87",x"c9",x"db"),
   588 => (x"ea",x"c2",x"1e",x"c0"),
   589 => (x"e2",x"fd",x"49",x"d4"),
   590 => (x"d0",x"ff",x"87",x"c2"),
   591 => (x"78",x"e0",x"c0",x"48"),
   592 => (x"1e",x"d4",x"ea",x"c2"),
   593 => (x"c1",x"4a",x"66",x"cc"),
   594 => (x"fc",x"c2",x"92",x"c8"),
   595 => (x"81",x"72",x"49",x"f0"),
   596 => (x"87",x"d2",x"c7",x"fe"),
   597 => (x"ac",x"c1",x"86",x"cc"),
   598 => (x"87",x"c4",x"c1",x"05"),
   599 => (x"c9",x"49",x"66",x"c4"),
   600 => (x"c4",x"1e",x"71",x"31"),
   601 => (x"c8",x"c1",x"4a",x"66"),
   602 => (x"f0",x"fc",x"c2",x"92"),
   603 => (x"fe",x"81",x"72",x"49"),
   604 => (x"c2",x"87",x"f9",x"ca"),
   605 => (x"c8",x"1e",x"d4",x"ea"),
   606 => (x"c8",x"c1",x"4a",x"66"),
   607 => (x"f0",x"fc",x"c2",x"92"),
   608 => (x"fe",x"81",x"72",x"49"),
   609 => (x"d7",x"87",x"d0",x"c5"),
   610 => (x"eb",x"d9",x"ff",x"49"),
   611 => (x"1e",x"c0",x"c8",x"87"),
   612 => (x"49",x"d4",x"ea",x"c2"),
   613 => (x"87",x"c1",x"e0",x"fd"),
   614 => (x"d0",x"ff",x"86",x"cc"),
   615 => (x"78",x"e0",x"c0",x"48"),
   616 => (x"4c",x"26",x"8e",x"f8"),
   617 => (x"4f",x"26",x"4b",x"26"),
   618 => (x"5c",x"5b",x"5e",x"0e"),
   619 => (x"86",x"fc",x"0e",x"5d"),
   620 => (x"d4",x"ff",x"4d",x"71"),
   621 => (x"7e",x"66",x"d4",x"4c"),
   622 => (x"a8",x"b7",x"c3",x"48"),
   623 => (x"87",x"e3",x"c1",x"01"),
   624 => (x"66",x"c4",x"1e",x"75"),
   625 => (x"93",x"c8",x"c1",x"4b"),
   626 => (x"83",x"f0",x"fc",x"c2"),
   627 => (x"fe",x"fd",x"49",x"73"),
   628 => (x"a3",x"c8",x"87",x"c7"),
   629 => (x"ff",x"49",x"69",x"49"),
   630 => (x"e1",x"c8",x"48",x"d0"),
   631 => (x"71",x"7c",x"dd",x"78"),
   632 => (x"98",x"ff",x"c3",x"48"),
   633 => (x"4a",x"71",x"7c",x"70"),
   634 => (x"72",x"2a",x"b7",x"c8"),
   635 => (x"98",x"ff",x"c3",x"48"),
   636 => (x"4a",x"71",x"7c",x"70"),
   637 => (x"72",x"2a",x"b7",x"d0"),
   638 => (x"98",x"ff",x"c3",x"48"),
   639 => (x"48",x"71",x"7c",x"70"),
   640 => (x"70",x"28",x"b7",x"d8"),
   641 => (x"7c",x"7c",x"c0",x"7c"),
   642 => (x"7c",x"7c",x"7c",x"7c"),
   643 => (x"7c",x"7c",x"7c",x"7c"),
   644 => (x"d0",x"ff",x"7c",x"7c"),
   645 => (x"78",x"e0",x"c0",x"48"),
   646 => (x"dc",x"1e",x"66",x"c4"),
   647 => (x"fc",x"d7",x"ff",x"49"),
   648 => (x"fc",x"86",x"c8",x"87"),
   649 => (x"26",x"4d",x"26",x"8e"),
   650 => (x"26",x"4b",x"26",x"4c"),
   651 => (x"1e",x"c0",x"1e",x"4f"),
   652 => (x"bf",x"c8",x"e9",x"c2"),
   653 => (x"87",x"f0",x"fd",x"49"),
   654 => (x"bf",x"cc",x"e9",x"c2"),
   655 => (x"e5",x"dc",x"fe",x"49"),
   656 => (x"fc",x"48",x"c0",x"87"),
   657 => (x"00",x"4f",x"26",x"8e"),
   658 => (x"00",x"00",x"2a",x"50"),
   659 => (x"00",x"00",x"2a",x"5c"),
   660 => (x"38",x"34",x"58",x"5a"),
   661 => (x"20",x"20",x"20",x"20"),
   662 => (x"00",x"44",x"48",x"56"),
   663 => (x"38",x"34",x"58",x"5a"),
   664 => (x"20",x"20",x"20",x"20"),
   665 => (x"00",x"4d",x"4f",x"52"),
   666 => (x"00",x"00",x"1d",x"8f"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

