
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom1 is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom1 is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"04",x"87",x"da",x"01"),
     1 => (x"58",x"0e",x"87",x"dd"),
     2 => (x"0e",x"5a",x"59",x"5e"),
     3 => (x"00",x"00",x"29",x"27"),
     4 => (x"4a",x"26",x"0f",x"00"),
     5 => (x"48",x"26",x"49",x"26"),
     6 => (x"08",x"26",x"80",x"ff"),
     7 => (x"00",x"2d",x"27",x"4f"),
     8 => (x"27",x"4f",x"00",x"00"),
     9 => (x"00",x"00",x"00",x"2a"),
    10 => (x"fd",x"00",x"4f",x"4f"),
    11 => (x"d0",x"c1",x"c3",x"87"),
    12 => (x"48",x"c0",x"c8",x"4e"),
    13 => (x"d5",x"c1",x"28",x"c2"),
    14 => (x"ea",x"d6",x"e5",x"ea"),
    15 => (x"c1",x"46",x"71",x"49"),
    16 => (x"87",x"f9",x"01",x"88"),
    17 => (x"49",x"d0",x"c1",x"c3"),
    18 => (x"48",x"ec",x"e9",x"c2"),
    19 => (x"03",x"89",x"d0",x"89"),
    20 => (x"40",x"40",x"40",x"c0"),
    21 => (x"d0",x"87",x"f6",x"40"),
    22 => (x"50",x"c0",x"05",x"81"),
    23 => (x"f9",x"05",x"89",x"c1"),
    24 => (x"ec",x"e9",x"c2",x"87"),
    25 => (x"e8",x"e9",x"c2",x"4d"),
    26 => (x"02",x"ad",x"74",x"4c"),
    27 => (x"0f",x"24",x"87",x"c4"),
    28 => (x"ef",x"c1",x"87",x"f7"),
    29 => (x"e9",x"c2",x"87",x"e6"),
    30 => (x"e9",x"c2",x"4d",x"ec"),
    31 => (x"ad",x"74",x"4c",x"ec"),
    32 => (x"c4",x"87",x"c6",x"02"),
    33 => (x"f5",x"0f",x"6c",x"8c"),
    34 => (x"87",x"fd",x"00",x"87"),
    35 => (x"71",x"86",x"fc",x"1e"),
    36 => (x"49",x"c0",x"ff",x"4a"),
    37 => (x"c0",x"c4",x"48",x"69"),
    38 => (x"48",x"7e",x"70",x"98"),
    39 => (x"87",x"f4",x"02",x"98"),
    40 => (x"fc",x"48",x"79",x"72"),
    41 => (x"0e",x"4f",x"26",x"8e"),
    42 => (x"0e",x"5c",x"5b",x"5e"),
    43 => (x"4c",x"c0",x"4b",x"71"),
    44 => (x"02",x"9a",x"4a",x"13"),
    45 => (x"49",x"72",x"87",x"cd"),
    46 => (x"c1",x"87",x"d1",x"ff"),
    47 => (x"9a",x"4a",x"13",x"84"),
    48 => (x"74",x"87",x"f3",x"05"),
    49 => (x"26",x"4c",x"26",x"48"),
    50 => (x"1e",x"4f",x"26",x"4b"),
    51 => (x"1e",x"73",x"1e",x"72"),
    52 => (x"02",x"11",x"48",x"12"),
    53 => (x"c3",x"4b",x"87",x"ca"),
    54 => (x"73",x"9b",x"98",x"df"),
    55 => (x"87",x"f0",x"02",x"88"),
    56 => (x"4a",x"26",x"4b",x"26"),
    57 => (x"73",x"1e",x"4f",x"26"),
    58 => (x"c1",x"1e",x"72",x"1e"),
    59 => (x"87",x"ca",x"04",x"8b"),
    60 => (x"02",x"11",x"48",x"12"),
    61 => (x"02",x"88",x"87",x"c4"),
    62 => (x"4a",x"26",x"87",x"f1"),
    63 => (x"4f",x"26",x"4b",x"26"),
    64 => (x"73",x"1e",x"74",x"1e"),
    65 => (x"c1",x"1e",x"72",x"1e"),
    66 => (x"87",x"d0",x"04",x"8b"),
    67 => (x"02",x"11",x"48",x"12"),
    68 => (x"c3",x"4c",x"87",x"ca"),
    69 => (x"74",x"9c",x"98",x"df"),
    70 => (x"87",x"eb",x"02",x"88"),
    71 => (x"4b",x"26",x"4a",x"26"),
    72 => (x"4f",x"26",x"4c",x"26"),
    73 => (x"81",x"48",x"73",x"1e"),
    74 => (x"c5",x"02",x"a9",x"73"),
    75 => (x"05",x"53",x"12",x"87"),
    76 => (x"4f",x"26",x"87",x"f6"),
    77 => (x"72",x"1e",x"73",x"1e"),
    78 => (x"e7",x"c0",x"02",x"9a"),
    79 => (x"c1",x"48",x"c0",x"87"),
    80 => (x"06",x"a9",x"72",x"4b"),
    81 => (x"82",x"72",x"87",x"d1"),
    82 => (x"73",x"87",x"c9",x"06"),
    83 => (x"01",x"a9",x"72",x"83"),
    84 => (x"87",x"c3",x"87",x"f4"),
    85 => (x"72",x"3a",x"b2",x"c1"),
    86 => (x"73",x"89",x"03",x"a9"),
    87 => (x"2a",x"c1",x"07",x"80"),
    88 => (x"87",x"f3",x"05",x"2b"),
    89 => (x"4f",x"26",x"4b",x"26"),
    90 => (x"c4",x"1e",x"75",x"1e"),
    91 => (x"a1",x"b7",x"71",x"4d"),
    92 => (x"c1",x"b9",x"ff",x"04"),
    93 => (x"07",x"bd",x"c3",x"81"),
    94 => (x"04",x"a2",x"b7",x"72"),
    95 => (x"82",x"c1",x"ba",x"ff"),
    96 => (x"fe",x"07",x"bd",x"c1"),
    97 => (x"2d",x"c1",x"87",x"ee"),
    98 => (x"c1",x"b8",x"ff",x"04"),
    99 => (x"04",x"2d",x"07",x"80"),
   100 => (x"81",x"c1",x"b9",x"ff"),
   101 => (x"26",x"4d",x"26",x"07"),
   102 => (x"1e",x"73",x"1e",x"4f"),
   103 => (x"66",x"c8",x"4a",x"71"),
   104 => (x"8b",x"c1",x"49",x"4b"),
   105 => (x"cf",x"02",x"99",x"71"),
   106 => (x"ff",x"48",x"12",x"87"),
   107 => (x"73",x"78",x"08",x"d4"),
   108 => (x"71",x"8b",x"c1",x"49"),
   109 => (x"87",x"f1",x"05",x"99"),
   110 => (x"4f",x"26",x"4b",x"26"),
   111 => (x"5c",x"5b",x"5e",x"0e"),
   112 => (x"ff",x"4a",x"71",x"0e"),
   113 => (x"66",x"cc",x"4c",x"d4"),
   114 => (x"8b",x"c1",x"49",x"4b"),
   115 => (x"ce",x"02",x"99",x"71"),
   116 => (x"7c",x"ff",x"c3",x"87"),
   117 => (x"49",x"73",x"52",x"6c"),
   118 => (x"99",x"71",x"8b",x"c1"),
   119 => (x"26",x"87",x"f2",x"05"),
   120 => (x"26",x"4b",x"26",x"4c"),
   121 => (x"1e",x"73",x"1e",x"4f"),
   122 => (x"c3",x"4b",x"d4",x"ff"),
   123 => (x"4a",x"6b",x"7b",x"ff"),
   124 => (x"6b",x"7b",x"ff",x"c3"),
   125 => (x"72",x"32",x"c8",x"49"),
   126 => (x"7b",x"ff",x"c3",x"b1"),
   127 => (x"31",x"c8",x"4a",x"6b"),
   128 => (x"ff",x"c3",x"b2",x"71"),
   129 => (x"c8",x"49",x"6b",x"7b"),
   130 => (x"71",x"b1",x"72",x"32"),
   131 => (x"26",x"4b",x"26",x"48"),
   132 => (x"5b",x"5e",x"0e",x"4f"),
   133 => (x"71",x"0e",x"5d",x"5c"),
   134 => (x"4c",x"d4",x"ff",x"4d"),
   135 => (x"ff",x"c3",x"48",x"75"),
   136 => (x"c2",x"7c",x"70",x"98"),
   137 => (x"05",x"bf",x"ec",x"e9"),
   138 => (x"66",x"d0",x"87",x"c8"),
   139 => (x"d4",x"30",x"c9",x"48"),
   140 => (x"66",x"d0",x"58",x"a6"),
   141 => (x"71",x"29",x"d8",x"49"),
   142 => (x"98",x"ff",x"c3",x"48"),
   143 => (x"66",x"d0",x"7c",x"70"),
   144 => (x"71",x"29",x"d0",x"49"),
   145 => (x"98",x"ff",x"c3",x"48"),
   146 => (x"66",x"d0",x"7c",x"70"),
   147 => (x"71",x"29",x"c8",x"49"),
   148 => (x"98",x"ff",x"c3",x"48"),
   149 => (x"66",x"d0",x"7c",x"70"),
   150 => (x"98",x"ff",x"c3",x"48"),
   151 => (x"49",x"75",x"7c",x"70"),
   152 => (x"48",x"71",x"29",x"d0"),
   153 => (x"70",x"98",x"ff",x"c3"),
   154 => (x"c9",x"4b",x"6c",x"7c"),
   155 => (x"c3",x"4a",x"ff",x"f0"),
   156 => (x"cf",x"05",x"ab",x"ff"),
   157 => (x"7c",x"71",x"49",x"87"),
   158 => (x"8a",x"c1",x"4b",x"6c"),
   159 => (x"71",x"87",x"c5",x"02"),
   160 => (x"87",x"f2",x"02",x"ab"),
   161 => (x"4d",x"26",x"48",x"73"),
   162 => (x"4b",x"26",x"4c",x"26"),
   163 => (x"c0",x"1e",x"4f",x"26"),
   164 => (x"48",x"d4",x"ff",x"49"),
   165 => (x"c1",x"78",x"ff",x"c3"),
   166 => (x"b7",x"c8",x"c3",x"81"),
   167 => (x"87",x"f1",x"04",x"a9"),
   168 => (x"5e",x"0e",x"4f",x"26"),
   169 => (x"0e",x"5d",x"5c",x"5b"),
   170 => (x"c1",x"f0",x"ff",x"c0"),
   171 => (x"c0",x"c1",x"4d",x"f7"),
   172 => (x"c0",x"c0",x"c0",x"c0"),
   173 => (x"87",x"d6",x"ff",x"4b"),
   174 => (x"4c",x"df",x"f8",x"c4"),
   175 => (x"49",x"75",x"1e",x"c0"),
   176 => (x"c4",x"87",x"ce",x"fd"),
   177 => (x"05",x"a8",x"c1",x"86"),
   178 => (x"ff",x"87",x"e5",x"c0"),
   179 => (x"ff",x"c3",x"48",x"d4"),
   180 => (x"c0",x"1e",x"73",x"78"),
   181 => (x"e9",x"c1",x"f0",x"e1"),
   182 => (x"87",x"f5",x"fc",x"49"),
   183 => (x"98",x"70",x"86",x"c4"),
   184 => (x"ff",x"87",x"ca",x"05"),
   185 => (x"ff",x"c3",x"48",x"d4"),
   186 => (x"cb",x"48",x"c1",x"78"),
   187 => (x"87",x"de",x"fe",x"87"),
   188 => (x"ff",x"05",x"8c",x"c1"),
   189 => (x"48",x"c0",x"87",x"c6"),
   190 => (x"4c",x"26",x"4d",x"26"),
   191 => (x"4f",x"26",x"4b",x"26"),
   192 => (x"5c",x"5b",x"5e",x"0e"),
   193 => (x"f0",x"ff",x"c0",x"0e"),
   194 => (x"ff",x"4c",x"c1",x"c1"),
   195 => (x"ff",x"c3",x"48",x"d4"),
   196 => (x"49",x"c4",x"cd",x"78"),
   197 => (x"d3",x"87",x"d0",x"f6"),
   198 => (x"74",x"1e",x"c0",x"4b"),
   199 => (x"87",x"f1",x"fb",x"49"),
   200 => (x"98",x"70",x"86",x"c4"),
   201 => (x"ff",x"87",x"ca",x"05"),
   202 => (x"ff",x"c3",x"48",x"d4"),
   203 => (x"cb",x"48",x"c1",x"78"),
   204 => (x"87",x"da",x"fd",x"87"),
   205 => (x"ff",x"05",x"8b",x"c1"),
   206 => (x"48",x"c0",x"87",x"df"),
   207 => (x"4b",x"26",x"4c",x"26"),
   208 => (x"00",x"00",x"4f",x"26"),
   209 => (x"00",x"44",x"4d",x"43"),
   210 => (x"5c",x"5b",x"5e",x"0e"),
   211 => (x"ff",x"c3",x"0e",x"5d"),
   212 => (x"4b",x"d4",x"ff",x"4d"),
   213 => (x"c6",x"87",x"f7",x"fc"),
   214 => (x"e1",x"c0",x"1e",x"ea"),
   215 => (x"49",x"c8",x"c1",x"f0"),
   216 => (x"c4",x"87",x"ee",x"fa"),
   217 => (x"02",x"a8",x"c1",x"86"),
   218 => (x"d3",x"fe",x"87",x"c8"),
   219 => (x"c1",x"48",x"c0",x"87"),
   220 => (x"f0",x"f9",x"87",x"e8"),
   221 => (x"cf",x"49",x"70",x"87"),
   222 => (x"c6",x"99",x"ff",x"ff"),
   223 => (x"c8",x"02",x"a9",x"ea"),
   224 => (x"87",x"fc",x"fd",x"87"),
   225 => (x"d1",x"c1",x"48",x"c0"),
   226 => (x"c0",x"7b",x"75",x"87"),
   227 => (x"d1",x"fc",x"4c",x"f1"),
   228 => (x"02",x"98",x"70",x"87"),
   229 => (x"c0",x"87",x"ec",x"c0"),
   230 => (x"f0",x"ff",x"c0",x"1e"),
   231 => (x"f9",x"49",x"fa",x"c1"),
   232 => (x"86",x"c4",x"87",x"ef"),
   233 => (x"da",x"05",x"98",x"70"),
   234 => (x"6b",x"7b",x"75",x"87"),
   235 => (x"75",x"7b",x"75",x"49"),
   236 => (x"75",x"7b",x"75",x"7b"),
   237 => (x"99",x"c0",x"c1",x"7b"),
   238 => (x"c1",x"87",x"c4",x"02"),
   239 => (x"c0",x"87",x"db",x"48"),
   240 => (x"c2",x"87",x"d7",x"48"),
   241 => (x"87",x"ca",x"05",x"ac"),
   242 => (x"f3",x"49",x"e4",x"cf"),
   243 => (x"48",x"c0",x"87",x"d9"),
   244 => (x"8c",x"c1",x"87",x"c8"),
   245 => (x"87",x"f6",x"fe",x"05"),
   246 => (x"4d",x"26",x"48",x"c0"),
   247 => (x"4b",x"26",x"4c",x"26"),
   248 => (x"00",x"00",x"4f",x"26"),
   249 => (x"43",x"48",x"44",x"53"),
   250 => (x"69",x"61",x"66",x"20"),
   251 => (x"00",x"0a",x"21",x"6c"),
   252 => (x"5c",x"5b",x"5e",x"0e"),
   253 => (x"d0",x"ff",x"0e",x"5d"),
   254 => (x"d0",x"e5",x"c0",x"4d"),
   255 => (x"c2",x"4c",x"c0",x"c1"),
   256 => (x"c1",x"48",x"ec",x"e9"),
   257 => (x"49",x"fc",x"d1",x"78"),
   258 => (x"c7",x"87",x"dc",x"f2"),
   259 => (x"f9",x"7d",x"c2",x"4b"),
   260 => (x"7d",x"c3",x"87",x"fc"),
   261 => (x"49",x"74",x"1e",x"c0"),
   262 => (x"c4",x"87",x"f6",x"f7"),
   263 => (x"05",x"a8",x"c1",x"86"),
   264 => (x"c2",x"4b",x"87",x"c1"),
   265 => (x"87",x"cb",x"05",x"ab"),
   266 => (x"f1",x"49",x"f4",x"d1"),
   267 => (x"48",x"c0",x"87",x"f9"),
   268 => (x"c1",x"87",x"f6",x"c0"),
   269 => (x"d4",x"ff",x"05",x"8b"),
   270 => (x"87",x"cc",x"fc",x"87"),
   271 => (x"58",x"f0",x"e9",x"c2"),
   272 => (x"cd",x"05",x"98",x"70"),
   273 => (x"c0",x"1e",x"c1",x"87"),
   274 => (x"d0",x"c1",x"f0",x"ff"),
   275 => (x"87",x"c1",x"f7",x"49"),
   276 => (x"d4",x"ff",x"86",x"c4"),
   277 => (x"78",x"ff",x"c3",x"48"),
   278 => (x"c2",x"87",x"cc",x"c5"),
   279 => (x"c2",x"58",x"f4",x"e9"),
   280 => (x"48",x"d4",x"ff",x"7d"),
   281 => (x"c1",x"78",x"ff",x"c3"),
   282 => (x"26",x"4d",x"26",x"48"),
   283 => (x"26",x"4b",x"26",x"4c"),
   284 => (x"00",x"00",x"00",x"4f"),
   285 => (x"52",x"52",x"45",x"49"),
   286 => (x"00",x"00",x"00",x"00"),
   287 => (x"00",x"49",x"50",x"53"),
   288 => (x"5c",x"5b",x"5e",x"0e"),
   289 => (x"4d",x"71",x"0e",x"5d"),
   290 => (x"ff",x"4c",x"ff",x"c3"),
   291 => (x"7b",x"74",x"4b",x"d4"),
   292 => (x"c4",x"48",x"d0",x"ff"),
   293 => (x"7b",x"74",x"78",x"c3"),
   294 => (x"ff",x"c0",x"1e",x"75"),
   295 => (x"49",x"d8",x"c1",x"f0"),
   296 => (x"c4",x"87",x"ee",x"f5"),
   297 => (x"02",x"98",x"70",x"86"),
   298 => (x"ec",x"d3",x"87",x"cb"),
   299 => (x"87",x"f7",x"ef",x"49"),
   300 => (x"ee",x"c0",x"48",x"c1"),
   301 => (x"c3",x"7b",x"74",x"87"),
   302 => (x"c0",x"c8",x"7b",x"fe"),
   303 => (x"49",x"66",x"d4",x"1e"),
   304 => (x"c4",x"87",x"d6",x"f3"),
   305 => (x"74",x"7b",x"74",x"86"),
   306 => (x"d8",x"7b",x"74",x"7b"),
   307 => (x"74",x"4a",x"e0",x"da"),
   308 => (x"c5",x"05",x"6b",x"7b"),
   309 => (x"05",x"8a",x"c1",x"87"),
   310 => (x"7b",x"74",x"87",x"f5"),
   311 => (x"c2",x"48",x"d0",x"ff"),
   312 => (x"26",x"48",x"c0",x"78"),
   313 => (x"26",x"4c",x"26",x"4d"),
   314 => (x"00",x"4f",x"26",x"4b"),
   315 => (x"74",x"69",x"72",x"57"),
   316 => (x"61",x"66",x"20",x"65"),
   317 => (x"64",x"65",x"6c",x"69"),
   318 => (x"5e",x"0e",x"00",x"0a"),
   319 => (x"0e",x"5d",x"5c",x"5b"),
   320 => (x"4b",x"71",x"86",x"fc"),
   321 => (x"c0",x"4c",x"d4",x"ff"),
   322 => (x"cd",x"ee",x"c5",x"7e"),
   323 => (x"ff",x"c3",x"4a",x"df"),
   324 => (x"c3",x"48",x"6c",x"7c"),
   325 => (x"c0",x"05",x"a8",x"fe"),
   326 => (x"4d",x"74",x"87",x"f8"),
   327 => (x"cc",x"02",x"9b",x"73"),
   328 => (x"1e",x"66",x"d4",x"87"),
   329 => (x"d3",x"f2",x"49",x"73"),
   330 => (x"d4",x"86",x"c4",x"87"),
   331 => (x"48",x"d0",x"ff",x"87"),
   332 => (x"d4",x"78",x"d1",x"c4"),
   333 => (x"ff",x"c3",x"4a",x"66"),
   334 => (x"05",x"8a",x"c1",x"7d"),
   335 => (x"a6",x"d8",x"87",x"f8"),
   336 => (x"7c",x"ff",x"c3",x"5a"),
   337 => (x"05",x"9b",x"73",x"7c"),
   338 => (x"d0",x"ff",x"87",x"c5"),
   339 => (x"c1",x"78",x"d0",x"48"),
   340 => (x"8a",x"c1",x"7e",x"4a"),
   341 => (x"87",x"f6",x"fe",x"05"),
   342 => (x"8e",x"fc",x"48",x"6e"),
   343 => (x"4c",x"26",x"4d",x"26"),
   344 => (x"4f",x"26",x"4b",x"26"),
   345 => (x"71",x"1e",x"73",x"1e"),
   346 => (x"ff",x"4b",x"c0",x"4a"),
   347 => (x"ff",x"c3",x"48",x"d4"),
   348 => (x"48",x"d0",x"ff",x"78"),
   349 => (x"ff",x"78",x"c3",x"c4"),
   350 => (x"ff",x"c3",x"48",x"d4"),
   351 => (x"c0",x"1e",x"72",x"78"),
   352 => (x"d1",x"c1",x"f0",x"ff"),
   353 => (x"87",x"c9",x"f2",x"49"),
   354 => (x"98",x"70",x"86",x"c4"),
   355 => (x"c8",x"87",x"d2",x"05"),
   356 => (x"66",x"cc",x"1e",x"c0"),
   357 => (x"87",x"e2",x"fd",x"49"),
   358 => (x"4b",x"70",x"86",x"c4"),
   359 => (x"c2",x"48",x"d0",x"ff"),
   360 => (x"26",x"48",x"73",x"78"),
   361 => (x"0e",x"4f",x"26",x"4b"),
   362 => (x"5d",x"5c",x"5b",x"5e"),
   363 => (x"c0",x"1e",x"c0",x"0e"),
   364 => (x"c9",x"c1",x"f0",x"ff"),
   365 => (x"87",x"d9",x"f1",x"49"),
   366 => (x"e9",x"c2",x"1e",x"d2"),
   367 => (x"f9",x"fc",x"49",x"f4"),
   368 => (x"c0",x"86",x"c8",x"87"),
   369 => (x"d2",x"84",x"c1",x"4c"),
   370 => (x"f8",x"04",x"ac",x"b7"),
   371 => (x"f4",x"e9",x"c2",x"87"),
   372 => (x"c3",x"49",x"bf",x"97"),
   373 => (x"c0",x"c1",x"99",x"c0"),
   374 => (x"e7",x"c0",x"05",x"a9"),
   375 => (x"fb",x"e9",x"c2",x"87"),
   376 => (x"d0",x"49",x"bf",x"97"),
   377 => (x"fc",x"e9",x"c2",x"31"),
   378 => (x"c8",x"4a",x"bf",x"97"),
   379 => (x"c2",x"b1",x"72",x"32"),
   380 => (x"bf",x"97",x"fd",x"e9"),
   381 => (x"4c",x"71",x"b1",x"4a"),
   382 => (x"ff",x"ff",x"ff",x"cf"),
   383 => (x"ca",x"84",x"c1",x"9c"),
   384 => (x"87",x"e7",x"c1",x"34"),
   385 => (x"97",x"fd",x"e9",x"c2"),
   386 => (x"31",x"c1",x"49",x"bf"),
   387 => (x"e9",x"c2",x"99",x"c6"),
   388 => (x"4a",x"bf",x"97",x"fe"),
   389 => (x"72",x"2a",x"b7",x"c7"),
   390 => (x"f9",x"e9",x"c2",x"b1"),
   391 => (x"4d",x"4a",x"bf",x"97"),
   392 => (x"e9",x"c2",x"9d",x"cf"),
   393 => (x"4a",x"bf",x"97",x"fa"),
   394 => (x"32",x"ca",x"9a",x"c3"),
   395 => (x"97",x"fb",x"e9",x"c2"),
   396 => (x"33",x"c2",x"4b",x"bf"),
   397 => (x"e9",x"c2",x"b2",x"73"),
   398 => (x"4b",x"bf",x"97",x"fc"),
   399 => (x"c6",x"9b",x"c0",x"c3"),
   400 => (x"b2",x"73",x"2b",x"b7"),
   401 => (x"48",x"c1",x"81",x"c2"),
   402 => (x"49",x"70",x"30",x"71"),
   403 => (x"30",x"75",x"48",x"c1"),
   404 => (x"4c",x"72",x"4d",x"70"),
   405 => (x"94",x"71",x"84",x"c1"),
   406 => (x"ad",x"b7",x"c0",x"c8"),
   407 => (x"c1",x"87",x"cc",x"06"),
   408 => (x"c8",x"2d",x"b7",x"34"),
   409 => (x"01",x"ad",x"b7",x"c0"),
   410 => (x"74",x"87",x"f4",x"ff"),
   411 => (x"26",x"4d",x"26",x"48"),
   412 => (x"26",x"4b",x"26",x"4c"),
   413 => (x"5b",x"5e",x"0e",x"4f"),
   414 => (x"f8",x"0e",x"5d",x"5c"),
   415 => (x"dc",x"f2",x"c2",x"86"),
   416 => (x"c2",x"78",x"c0",x"48"),
   417 => (x"c0",x"1e",x"d4",x"ea"),
   418 => (x"87",x"d8",x"fb",x"49"),
   419 => (x"98",x"70",x"86",x"c4"),
   420 => (x"c0",x"87",x"c5",x"05"),
   421 => (x"87",x"c0",x"c9",x"48"),
   422 => (x"7e",x"c1",x"4d",x"c0"),
   423 => (x"bf",x"f8",x"fe",x"c0"),
   424 => (x"ca",x"eb",x"c2",x"49"),
   425 => (x"4b",x"c8",x"71",x"4a"),
   426 => (x"70",x"87",x"fb",x"e8"),
   427 => (x"87",x"c2",x"05",x"98"),
   428 => (x"fe",x"c0",x"7e",x"c0"),
   429 => (x"c2",x"49",x"bf",x"f4"),
   430 => (x"71",x"4a",x"e6",x"eb"),
   431 => (x"e5",x"e8",x"4b",x"c8"),
   432 => (x"05",x"98",x"70",x"87"),
   433 => (x"7e",x"c0",x"87",x"c2"),
   434 => (x"fd",x"c0",x"02",x"6e"),
   435 => (x"da",x"f1",x"c2",x"87"),
   436 => (x"f2",x"c2",x"4d",x"bf"),
   437 => (x"7e",x"bf",x"9f",x"d2"),
   438 => (x"ea",x"d6",x"c5",x"48"),
   439 => (x"87",x"c7",x"05",x"a8"),
   440 => (x"bf",x"da",x"f1",x"c2"),
   441 => (x"6e",x"87",x"ce",x"4d"),
   442 => (x"d5",x"e9",x"ca",x"48"),
   443 => (x"87",x"c5",x"02",x"a8"),
   444 => (x"e3",x"c7",x"48",x"c0"),
   445 => (x"d4",x"ea",x"c2",x"87"),
   446 => (x"f9",x"49",x"75",x"1e"),
   447 => (x"86",x"c4",x"87",x"e6"),
   448 => (x"c5",x"05",x"98",x"70"),
   449 => (x"c7",x"48",x"c0",x"87"),
   450 => (x"fe",x"c0",x"87",x"ce"),
   451 => (x"c2",x"49",x"bf",x"f4"),
   452 => (x"71",x"4a",x"e6",x"eb"),
   453 => (x"cd",x"e7",x"4b",x"c8"),
   454 => (x"05",x"98",x"70",x"87"),
   455 => (x"f2",x"c2",x"87",x"c8"),
   456 => (x"78",x"c1",x"48",x"dc"),
   457 => (x"fe",x"c0",x"87",x"da"),
   458 => (x"c2",x"49",x"bf",x"f8"),
   459 => (x"71",x"4a",x"ca",x"eb"),
   460 => (x"f1",x"e6",x"4b",x"c8"),
   461 => (x"02",x"98",x"70",x"87"),
   462 => (x"c0",x"87",x"c5",x"c0"),
   463 => (x"87",x"d8",x"c6",x"48"),
   464 => (x"97",x"d2",x"f2",x"c2"),
   465 => (x"d5",x"c1",x"49",x"bf"),
   466 => (x"cd",x"c0",x"05",x"a9"),
   467 => (x"d3",x"f2",x"c2",x"87"),
   468 => (x"c2",x"49",x"bf",x"97"),
   469 => (x"c0",x"02",x"a9",x"ea"),
   470 => (x"48",x"c0",x"87",x"c5"),
   471 => (x"c2",x"87",x"f9",x"c5"),
   472 => (x"bf",x"97",x"d4",x"ea"),
   473 => (x"e9",x"c3",x"48",x"7e"),
   474 => (x"ce",x"c0",x"02",x"a8"),
   475 => (x"c3",x"48",x"6e",x"87"),
   476 => (x"c0",x"02",x"a8",x"eb"),
   477 => (x"48",x"c0",x"87",x"c5"),
   478 => (x"c2",x"87",x"dd",x"c5"),
   479 => (x"bf",x"97",x"df",x"ea"),
   480 => (x"c0",x"05",x"99",x"49"),
   481 => (x"ea",x"c2",x"87",x"cc"),
   482 => (x"49",x"bf",x"97",x"e0"),
   483 => (x"c0",x"02",x"a9",x"c2"),
   484 => (x"48",x"c0",x"87",x"c5"),
   485 => (x"c2",x"87",x"c1",x"c5"),
   486 => (x"bf",x"97",x"e1",x"ea"),
   487 => (x"d8",x"f2",x"c2",x"48"),
   488 => (x"48",x"4c",x"70",x"58"),
   489 => (x"f2",x"c2",x"88",x"c1"),
   490 => (x"ea",x"c2",x"58",x"dc"),
   491 => (x"49",x"bf",x"97",x"e2"),
   492 => (x"ea",x"c2",x"81",x"75"),
   493 => (x"4a",x"bf",x"97",x"e3"),
   494 => (x"a1",x"72",x"32",x"c8"),
   495 => (x"ec",x"f6",x"c2",x"7e"),
   496 => (x"c2",x"78",x"6e",x"48"),
   497 => (x"bf",x"97",x"e4",x"ea"),
   498 => (x"58",x"a6",x"c8",x"48"),
   499 => (x"bf",x"dc",x"f2",x"c2"),
   500 => (x"87",x"cf",x"c2",x"02"),
   501 => (x"bf",x"f4",x"fe",x"c0"),
   502 => (x"e6",x"eb",x"c2",x"49"),
   503 => (x"4b",x"c8",x"71",x"4a"),
   504 => (x"70",x"87",x"c3",x"e4"),
   505 => (x"c5",x"c0",x"02",x"98"),
   506 => (x"c3",x"48",x"c0",x"87"),
   507 => (x"f2",x"c2",x"87",x"ea"),
   508 => (x"c2",x"4c",x"bf",x"d4"),
   509 => (x"c2",x"5c",x"c0",x"f7"),
   510 => (x"bf",x"97",x"f9",x"ea"),
   511 => (x"c2",x"31",x"c8",x"49"),
   512 => (x"bf",x"97",x"f8",x"ea"),
   513 => (x"c2",x"49",x"a1",x"4a"),
   514 => (x"bf",x"97",x"fa",x"ea"),
   515 => (x"72",x"32",x"d0",x"4a"),
   516 => (x"ea",x"c2",x"49",x"a1"),
   517 => (x"4a",x"bf",x"97",x"fb"),
   518 => (x"a1",x"72",x"32",x"d8"),
   519 => (x"91",x"66",x"c4",x"49"),
   520 => (x"bf",x"ec",x"f6",x"c2"),
   521 => (x"f4",x"f6",x"c2",x"81"),
   522 => (x"c1",x"eb",x"c2",x"59"),
   523 => (x"c8",x"4a",x"bf",x"97"),
   524 => (x"c0",x"eb",x"c2",x"32"),
   525 => (x"a2",x"4b",x"bf",x"97"),
   526 => (x"c2",x"eb",x"c2",x"4a"),
   527 => (x"d0",x"4b",x"bf",x"97"),
   528 => (x"4a",x"a2",x"73",x"33"),
   529 => (x"97",x"c3",x"eb",x"c2"),
   530 => (x"9b",x"cf",x"4b",x"bf"),
   531 => (x"a2",x"73",x"33",x"d8"),
   532 => (x"f8",x"f6",x"c2",x"4a"),
   533 => (x"74",x"8a",x"c2",x"5a"),
   534 => (x"f8",x"f6",x"c2",x"92"),
   535 => (x"78",x"a1",x"72",x"48"),
   536 => (x"c2",x"87",x"c1",x"c1"),
   537 => (x"bf",x"97",x"e6",x"ea"),
   538 => (x"c2",x"31",x"c8",x"49"),
   539 => (x"bf",x"97",x"e5",x"ea"),
   540 => (x"c5",x"49",x"a1",x"4a"),
   541 => (x"81",x"ff",x"c7",x"31"),
   542 => (x"f7",x"c2",x"29",x"c9"),
   543 => (x"ea",x"c2",x"59",x"c0"),
   544 => (x"4a",x"bf",x"97",x"eb"),
   545 => (x"ea",x"c2",x"32",x"c8"),
   546 => (x"4b",x"bf",x"97",x"ea"),
   547 => (x"66",x"c4",x"4a",x"a2"),
   548 => (x"c2",x"82",x"6e",x"92"),
   549 => (x"c2",x"5a",x"fc",x"f6"),
   550 => (x"c0",x"48",x"f4",x"f6"),
   551 => (x"f0",x"f6",x"c2",x"78"),
   552 => (x"78",x"a1",x"72",x"48"),
   553 => (x"48",x"c0",x"f7",x"c2"),
   554 => (x"bf",x"f4",x"f6",x"c2"),
   555 => (x"c4",x"f7",x"c2",x"78"),
   556 => (x"f8",x"f6",x"c2",x"48"),
   557 => (x"f2",x"c2",x"78",x"bf"),
   558 => (x"c0",x"02",x"bf",x"dc"),
   559 => (x"48",x"74",x"87",x"c9"),
   560 => (x"7e",x"70",x"30",x"c4"),
   561 => (x"c2",x"87",x"c9",x"c0"),
   562 => (x"48",x"bf",x"fc",x"f6"),
   563 => (x"7e",x"70",x"30",x"c4"),
   564 => (x"48",x"e0",x"f2",x"c2"),
   565 => (x"48",x"c1",x"78",x"6e"),
   566 => (x"4d",x"26",x"8e",x"f8"),
   567 => (x"4b",x"26",x"4c",x"26"),
   568 => (x"5e",x"0e",x"4f",x"26"),
   569 => (x"0e",x"5d",x"5c",x"5b"),
   570 => (x"f2",x"c2",x"4a",x"71"),
   571 => (x"cb",x"02",x"bf",x"dc"),
   572 => (x"c7",x"4b",x"72",x"87"),
   573 => (x"c1",x"4d",x"72",x"2b"),
   574 => (x"87",x"c9",x"9d",x"ff"),
   575 => (x"2b",x"c8",x"4b",x"72"),
   576 => (x"ff",x"c3",x"4d",x"72"),
   577 => (x"ec",x"f6",x"c2",x"9d"),
   578 => (x"fe",x"c0",x"83",x"bf"),
   579 => (x"02",x"ab",x"bf",x"f0"),
   580 => (x"fe",x"c0",x"87",x"d9"),
   581 => (x"ea",x"c2",x"5b",x"f4"),
   582 => (x"49",x"73",x"1e",x"d4"),
   583 => (x"c4",x"87",x"c5",x"f1"),
   584 => (x"05",x"98",x"70",x"86"),
   585 => (x"48",x"c0",x"87",x"c5"),
   586 => (x"c2",x"87",x"e6",x"c0"),
   587 => (x"02",x"bf",x"dc",x"f2"),
   588 => (x"49",x"75",x"87",x"d2"),
   589 => (x"ea",x"c2",x"91",x"c4"),
   590 => (x"4c",x"69",x"81",x"d4"),
   591 => (x"ff",x"ff",x"ff",x"cf"),
   592 => (x"87",x"cb",x"9c",x"ff"),
   593 => (x"91",x"c2",x"49",x"75"),
   594 => (x"81",x"d4",x"ea",x"c2"),
   595 => (x"74",x"4c",x"69",x"9f"),
   596 => (x"26",x"4d",x"26",x"48"),
   597 => (x"26",x"4b",x"26",x"4c"),
   598 => (x"5b",x"5e",x"0e",x"4f"),
   599 => (x"f0",x"0e",x"5d",x"5c"),
   600 => (x"59",x"a6",x"cc",x"86"),
   601 => (x"c5",x"05",x"66",x"c8"),
   602 => (x"c4",x"48",x"c0",x"87"),
   603 => (x"66",x"c8",x"87",x"c4"),
   604 => (x"70",x"80",x"c8",x"48"),
   605 => (x"78",x"c0",x"48",x"7e"),
   606 => (x"02",x"66",x"e0",x"c0"),
   607 => (x"e0",x"c0",x"87",x"c8"),
   608 => (x"05",x"bf",x"97",x"66"),
   609 => (x"48",x"c0",x"87",x"c5"),
   610 => (x"c0",x"87",x"e7",x"c3"),
   611 => (x"49",x"49",x"c1",x"1e"),
   612 => (x"c4",x"87",x"e5",x"d0"),
   613 => (x"9c",x"4c",x"70",x"86"),
   614 => (x"87",x"fe",x"c0",x"02"),
   615 => (x"4a",x"e4",x"f2",x"c2"),
   616 => (x"49",x"66",x"e0",x"c0"),
   617 => (x"87",x"e3",x"dc",x"ff"),
   618 => (x"c0",x"02",x"98",x"70"),
   619 => (x"4a",x"74",x"87",x"ec"),
   620 => (x"49",x"66",x"e0",x"c0"),
   621 => (x"dd",x"ff",x"4b",x"cb"),
   622 => (x"98",x"70",x"87",x"c6"),
   623 => (x"c0",x"87",x"db",x"02"),
   624 => (x"02",x"9c",x"74",x"1e"),
   625 => (x"4d",x"c0",x"87",x"c4"),
   626 => (x"4d",x"c1",x"87",x"c2"),
   627 => (x"e7",x"cf",x"49",x"75"),
   628 => (x"70",x"86",x"c4",x"87"),
   629 => (x"ff",x"05",x"9c",x"4c"),
   630 => (x"9c",x"74",x"87",x"c2"),
   631 => (x"87",x"d0",x"c2",x"02"),
   632 => (x"6e",x"49",x"a4",x"dc"),
   633 => (x"da",x"78",x"69",x"48"),
   634 => (x"66",x"c8",x"49",x"a4"),
   635 => (x"c8",x"80",x"c4",x"48"),
   636 => (x"69",x"9f",x"58",x"a6"),
   637 => (x"08",x"66",x"c4",x"48"),
   638 => (x"dc",x"f2",x"c2",x"78"),
   639 => (x"87",x"d2",x"02",x"bf"),
   640 => (x"9f",x"49",x"a4",x"d4"),
   641 => (x"ff",x"c0",x"49",x"69"),
   642 => (x"48",x"71",x"99",x"ff"),
   643 => (x"58",x"a6",x"30",x"d0"),
   644 => (x"a6",x"cc",x"87",x"c5"),
   645 => (x"cc",x"78",x"c0",x"48"),
   646 => (x"66",x"c4",x"48",x"66"),
   647 => (x"66",x"c4",x"80",x"bf"),
   648 => (x"66",x"c8",x"78",x"08"),
   649 => (x"c8",x"78",x"c0",x"48"),
   650 => (x"81",x"cc",x"49",x"66"),
   651 => (x"79",x"bf",x"66",x"c4"),
   652 => (x"d0",x"49",x"66",x"c8"),
   653 => (x"4d",x"79",x"c0",x"81"),
   654 => (x"c8",x"4c",x"66",x"c4"),
   655 => (x"82",x"d4",x"4a",x"66"),
   656 => (x"91",x"c8",x"49",x"75"),
   657 => (x"c0",x"49",x"a1",x"72"),
   658 => (x"c1",x"79",x"6c",x"41"),
   659 => (x"ad",x"b7",x"c6",x"85"),
   660 => (x"87",x"e7",x"ff",x"04"),
   661 => (x"c9",x"4a",x"bf",x"6e"),
   662 => (x"c0",x"49",x"72",x"2a"),
   663 => (x"db",x"ff",x"4a",x"f0"),
   664 => (x"4a",x"70",x"87",x"d2"),
   665 => (x"c1",x"49",x"66",x"c8"),
   666 => (x"79",x"72",x"81",x"c4"),
   667 => (x"87",x"c2",x"48",x"c1"),
   668 => (x"8e",x"f0",x"48",x"c0"),
   669 => (x"4c",x"26",x"4d",x"26"),
   670 => (x"4f",x"26",x"4b",x"26"),
   671 => (x"5c",x"5b",x"5e",x"0e"),
   672 => (x"4c",x"71",x"0e",x"5d"),
   673 => (x"74",x"4d",x"66",x"d0"),
   674 => (x"c2",x"c1",x"02",x"9c"),
   675 => (x"49",x"a4",x"c8",x"87"),
   676 => (x"fa",x"c0",x"02",x"69"),
   677 => (x"85",x"49",x"6c",x"87"),
   678 => (x"f2",x"c2",x"b9",x"75"),
   679 => (x"ff",x"4a",x"bf",x"d8"),
   680 => (x"71",x"99",x"72",x"ba"),
   681 => (x"e4",x"c0",x"02",x"99"),
   682 => (x"4b",x"a4",x"c4",x"87"),
   683 => (x"f1",x"f8",x"49",x"6b"),
   684 => (x"c2",x"7b",x"70",x"87"),
   685 => (x"49",x"bf",x"d4",x"f2"),
   686 => (x"7c",x"71",x"81",x"6c"),
   687 => (x"f2",x"c2",x"b9",x"75"),
   688 => (x"ff",x"4a",x"bf",x"d8"),
   689 => (x"71",x"99",x"72",x"ba"),
   690 => (x"dc",x"ff",x"05",x"99"),
   691 => (x"26",x"7c",x"75",x"87"),
   692 => (x"26",x"4c",x"26",x"4d"),
   693 => (x"1e",x"4f",x"26",x"4b"),
   694 => (x"4b",x"71",x"1e",x"73"),
   695 => (x"87",x"c7",x"02",x"9b"),
   696 => (x"69",x"49",x"a3",x"c8"),
   697 => (x"c0",x"87",x"c5",x"05"),
   698 => (x"87",x"f6",x"c0",x"48"),
   699 => (x"bf",x"f0",x"f6",x"c2"),
   700 => (x"4a",x"a3",x"c4",x"49"),
   701 => (x"8a",x"c2",x"4a",x"6a"),
   702 => (x"bf",x"d4",x"f2",x"c2"),
   703 => (x"49",x"a1",x"72",x"92"),
   704 => (x"bf",x"d8",x"f2",x"c2"),
   705 => (x"72",x"9a",x"6b",x"4a"),
   706 => (x"fe",x"c0",x"49",x"a1"),
   707 => (x"66",x"c8",x"59",x"f4"),
   708 => (x"cf",x"e9",x"71",x"1e"),
   709 => (x"70",x"86",x"c4",x"87"),
   710 => (x"87",x"c4",x"05",x"98"),
   711 => (x"87",x"c2",x"48",x"c0"),
   712 => (x"4b",x"26",x"48",x"c1"),
   713 => (x"73",x"1e",x"4f",x"26"),
   714 => (x"9b",x"4b",x"71",x"1e"),
   715 => (x"c8",x"87",x"c7",x"02"),
   716 => (x"05",x"69",x"49",x"a3"),
   717 => (x"48",x"c0",x"87",x"c5"),
   718 => (x"c2",x"87",x"f6",x"c0"),
   719 => (x"49",x"bf",x"f0",x"f6"),
   720 => (x"6a",x"4a",x"a3",x"c4"),
   721 => (x"c2",x"8a",x"c2",x"4a"),
   722 => (x"92",x"bf",x"d4",x"f2"),
   723 => (x"c2",x"49",x"a1",x"72"),
   724 => (x"4a",x"bf",x"d8",x"f2"),
   725 => (x"a1",x"72",x"9a",x"6b"),
   726 => (x"f4",x"fe",x"c0",x"49"),
   727 => (x"1e",x"66",x"c8",x"59"),
   728 => (x"87",x"dc",x"e4",x"71"),
   729 => (x"98",x"70",x"86",x"c4"),
   730 => (x"c0",x"87",x"c4",x"05"),
   731 => (x"c1",x"87",x"c2",x"48"),
   732 => (x"26",x"4b",x"26",x"48"),
   733 => (x"5b",x"5e",x"0e",x"4f"),
   734 => (x"f8",x"0e",x"5d",x"5c"),
   735 => (x"c4",x"7e",x"71",x"86"),
   736 => (x"78",x"ff",x"48",x"a6"),
   737 => (x"ff",x"ff",x"ff",x"c1"),
   738 => (x"c0",x"4d",x"ff",x"ff"),
   739 => (x"d4",x"4a",x"6e",x"4b"),
   740 => (x"c8",x"49",x"73",x"82"),
   741 => (x"49",x"a1",x"72",x"91"),
   742 => (x"69",x"4c",x"66",x"d8"),
   743 => (x"ac",x"b7",x"c0",x"8c"),
   744 => (x"75",x"87",x"cb",x"04"),
   745 => (x"c5",x"03",x"ac",x"b7"),
   746 => (x"5b",x"a6",x"c8",x"87"),
   747 => (x"83",x"c1",x"4d",x"74"),
   748 => (x"04",x"ab",x"b7",x"c6"),
   749 => (x"c4",x"87",x"d6",x"ff"),
   750 => (x"8e",x"f8",x"48",x"66"),
   751 => (x"4c",x"26",x"4d",x"26"),
   752 => (x"4f",x"26",x"4b",x"26"),
   753 => (x"5c",x"5b",x"5e",x"0e"),
   754 => (x"86",x"f0",x"0e",x"5d"),
   755 => (x"a6",x"c4",x"7e",x"71"),
   756 => (x"ff",x"ff",x"c1",x"48"),
   757 => (x"78",x"ff",x"ff",x"ff"),
   758 => (x"78",x"ff",x"80",x"c4"),
   759 => (x"4c",x"c0",x"4d",x"c0"),
   760 => (x"83",x"d4",x"4b",x"6e"),
   761 => (x"92",x"c8",x"4a",x"74"),
   762 => (x"75",x"4a",x"a2",x"73"),
   763 => (x"73",x"91",x"c8",x"49"),
   764 => (x"48",x"6a",x"49",x"a1"),
   765 => (x"a6",x"d0",x"88",x"69"),
   766 => (x"02",x"ad",x"74",x"58"),
   767 => (x"66",x"c4",x"87",x"cf"),
   768 => (x"87",x"c9",x"03",x"a8"),
   769 => (x"c4",x"5c",x"a6",x"cc"),
   770 => (x"66",x"cc",x"48",x"a6"),
   771 => (x"c6",x"84",x"c1",x"78"),
   772 => (x"ff",x"04",x"ac",x"b7"),
   773 => (x"85",x"c1",x"87",x"ca"),
   774 => (x"04",x"ad",x"b7",x"c6"),
   775 => (x"c8",x"87",x"ff",x"fe"),
   776 => (x"8e",x"f0",x"48",x"66"),
   777 => (x"4c",x"26",x"4d",x"26"),
   778 => (x"4f",x"26",x"4b",x"26"),
   779 => (x"5c",x"5b",x"5e",x"0e"),
   780 => (x"86",x"ec",x"0e",x"5d"),
   781 => (x"e4",x"c0",x"4b",x"71"),
   782 => (x"28",x"c9",x"48",x"66"),
   783 => (x"c2",x"58",x"a6",x"c8"),
   784 => (x"4a",x"bf",x"d8",x"f2"),
   785 => (x"48",x"72",x"ba",x"ff"),
   786 => (x"cc",x"98",x"66",x"c4"),
   787 => (x"9b",x"73",x"58",x"a6"),
   788 => (x"87",x"c1",x"c3",x"02"),
   789 => (x"69",x"49",x"a3",x"c8"),
   790 => (x"87",x"f9",x"c2",x"02"),
   791 => (x"98",x"6b",x"48",x"72"),
   792 => (x"c4",x"58",x"a6",x"d4"),
   793 => (x"7e",x"6c",x"4c",x"a3"),
   794 => (x"d0",x"48",x"66",x"c8"),
   795 => (x"c6",x"05",x"a8",x"66"),
   796 => (x"7b",x"66",x"c4",x"87"),
   797 => (x"c8",x"87",x"cc",x"c2"),
   798 => (x"49",x"73",x"1e",x"66"),
   799 => (x"c4",x"87",x"f6",x"fb"),
   800 => (x"c0",x"4d",x"70",x"86"),
   801 => (x"d0",x"04",x"ad",x"b7"),
   802 => (x"4a",x"a3",x"d4",x"87"),
   803 => (x"91",x"c8",x"49",x"75"),
   804 => (x"21",x"49",x"a1",x"72"),
   805 => (x"c7",x"7c",x"69",x"7b"),
   806 => (x"cc",x"7b",x"c0",x"87"),
   807 => (x"7c",x"69",x"49",x"a3"),
   808 => (x"6b",x"48",x"66",x"c4"),
   809 => (x"58",x"a6",x"c8",x"88"),
   810 => (x"73",x"1e",x"66",x"d0"),
   811 => (x"87",x"c5",x"fb",x"49"),
   812 => (x"4d",x"70",x"86",x"c4"),
   813 => (x"49",x"a3",x"c4",x"c1"),
   814 => (x"69",x"48",x"a6",x"c8"),
   815 => (x"48",x"66",x"d0",x"78"),
   816 => (x"06",x"a8",x"66",x"c8"),
   817 => (x"c0",x"87",x"f2",x"c0"),
   818 => (x"c0",x"04",x"ad",x"b7"),
   819 => (x"a6",x"cc",x"87",x"eb"),
   820 => (x"78",x"a3",x"d4",x"48"),
   821 => (x"91",x"c8",x"49",x"75"),
   822 => (x"d0",x"81",x"66",x"cc"),
   823 => (x"88",x"69",x"48",x"66"),
   824 => (x"66",x"c8",x"49",x"70"),
   825 => (x"87",x"d1",x"06",x"a9"),
   826 => (x"d7",x"fb",x"49",x"73"),
   827 => (x"c8",x"49",x"70",x"87"),
   828 => (x"81",x"66",x"cc",x"91"),
   829 => (x"6e",x"41",x"66",x"d0"),
   830 => (x"1e",x"66",x"c4",x"79"),
   831 => (x"fb",x"f5",x"49",x"73"),
   832 => (x"c2",x"86",x"c4",x"87"),
   833 => (x"73",x"1e",x"d4",x"ea"),
   834 => (x"87",x"cb",x"f7",x"49"),
   835 => (x"a3",x"d0",x"86",x"c4"),
   836 => (x"66",x"e4",x"c0",x"49"),
   837 => (x"26",x"8e",x"ec",x"79"),
   838 => (x"26",x"4c",x"26",x"4d"),
   839 => (x"1e",x"4f",x"26",x"4b"),
   840 => (x"4b",x"71",x"1e",x"73"),
   841 => (x"e4",x"c0",x"02",x"9b"),
   842 => (x"c4",x"f7",x"c2",x"87"),
   843 => (x"c2",x"4a",x"73",x"5b"),
   844 => (x"d4",x"f2",x"c2",x"8a"),
   845 => (x"c2",x"92",x"49",x"bf"),
   846 => (x"48",x"bf",x"f0",x"f6"),
   847 => (x"f7",x"c2",x"80",x"72"),
   848 => (x"48",x"71",x"58",x"c8"),
   849 => (x"f2",x"c2",x"30",x"c4"),
   850 => (x"ed",x"c0",x"58",x"e4"),
   851 => (x"c0",x"f7",x"c2",x"87"),
   852 => (x"f4",x"f6",x"c2",x"48"),
   853 => (x"f7",x"c2",x"78",x"bf"),
   854 => (x"f6",x"c2",x"48",x"c4"),
   855 => (x"c2",x"78",x"bf",x"f8"),
   856 => (x"02",x"bf",x"dc",x"f2"),
   857 => (x"f2",x"c2",x"87",x"c9"),
   858 => (x"c4",x"49",x"bf",x"d4"),
   859 => (x"c2",x"87",x"c7",x"31"),
   860 => (x"49",x"bf",x"fc",x"f6"),
   861 => (x"f2",x"c2",x"31",x"c4"),
   862 => (x"4b",x"26",x"59",x"e4"),
   863 => (x"5e",x"0e",x"4f",x"26"),
   864 => (x"71",x"0e",x"5c",x"5b"),
   865 => (x"72",x"4b",x"c0",x"4a"),
   866 => (x"e0",x"c0",x"02",x"9a"),
   867 => (x"49",x"a2",x"da",x"87"),
   868 => (x"c2",x"4b",x"69",x"9f"),
   869 => (x"02",x"bf",x"dc",x"f2"),
   870 => (x"a2",x"d4",x"87",x"cf"),
   871 => (x"49",x"69",x"9f",x"49"),
   872 => (x"ff",x"ff",x"c0",x"4c"),
   873 => (x"c2",x"34",x"d0",x"9c"),
   874 => (x"74",x"4c",x"c0",x"87"),
   875 => (x"fd",x"49",x"73",x"b3"),
   876 => (x"4c",x"26",x"87",x"ed"),
   877 => (x"4f",x"26",x"4b",x"26"),
   878 => (x"5c",x"5b",x"5e",x"0e"),
   879 => (x"86",x"f0",x"0e",x"5d"),
   880 => (x"cf",x"59",x"a6",x"c8"),
   881 => (x"f8",x"ff",x"ff",x"ff"),
   882 => (x"c4",x"7e",x"c0",x"4c"),
   883 => (x"87",x"d8",x"02",x"66"),
   884 => (x"48",x"d0",x"ea",x"c2"),
   885 => (x"ea",x"c2",x"78",x"c0"),
   886 => (x"f7",x"c2",x"48",x"c8"),
   887 => (x"c2",x"78",x"bf",x"c4"),
   888 => (x"c2",x"48",x"cc",x"ea"),
   889 => (x"78",x"bf",x"c0",x"f7"),
   890 => (x"48",x"f1",x"f2",x"c2"),
   891 => (x"f2",x"c2",x"50",x"c0"),
   892 => (x"c2",x"49",x"bf",x"e0"),
   893 => (x"4a",x"bf",x"d0",x"ea"),
   894 => (x"c4",x"03",x"aa",x"71"),
   895 => (x"49",x"72",x"87",x"cc"),
   896 => (x"c0",x"05",x"99",x"cf"),
   897 => (x"fe",x"c0",x"87",x"ea"),
   898 => (x"ea",x"c2",x"48",x"f0"),
   899 => (x"c2",x"78",x"bf",x"c8"),
   900 => (x"c2",x"1e",x"d4",x"ea"),
   901 => (x"49",x"bf",x"c8",x"ea"),
   902 => (x"48",x"c8",x"ea",x"c2"),
   903 => (x"71",x"78",x"a1",x"c1"),
   904 => (x"87",x"c0",x"dd",x"ff"),
   905 => (x"fe",x"c0",x"86",x"c4"),
   906 => (x"ea",x"c2",x"48",x"ec"),
   907 => (x"87",x"cc",x"78",x"d4"),
   908 => (x"bf",x"ec",x"fe",x"c0"),
   909 => (x"80",x"e0",x"c0",x"48"),
   910 => (x"58",x"f0",x"fe",x"c0"),
   911 => (x"bf",x"d0",x"ea",x"c2"),
   912 => (x"c2",x"80",x"c1",x"48"),
   913 => (x"27",x"58",x"d4",x"ea"),
   914 => (x"00",x"00",x"0f",x"ac"),
   915 => (x"4d",x"bf",x"97",x"bf"),
   916 => (x"e5",x"c2",x"02",x"9d"),
   917 => (x"ad",x"e5",x"c3",x"87"),
   918 => (x"87",x"de",x"c2",x"02"),
   919 => (x"bf",x"ec",x"fe",x"c0"),
   920 => (x"49",x"a3",x"cb",x"4b"),
   921 => (x"ac",x"cf",x"4c",x"11"),
   922 => (x"87",x"d2",x"c1",x"05"),
   923 => (x"99",x"df",x"49",x"75"),
   924 => (x"91",x"cd",x"89",x"c1"),
   925 => (x"81",x"e4",x"f2",x"c2"),
   926 => (x"12",x"4a",x"a3",x"c1"),
   927 => (x"4a",x"a3",x"c3",x"51"),
   928 => (x"a3",x"c5",x"51",x"12"),
   929 => (x"c7",x"51",x"12",x"4a"),
   930 => (x"51",x"12",x"4a",x"a3"),
   931 => (x"12",x"4a",x"a3",x"c9"),
   932 => (x"4a",x"a3",x"ce",x"51"),
   933 => (x"a3",x"d0",x"51",x"12"),
   934 => (x"d2",x"51",x"12",x"4a"),
   935 => (x"51",x"12",x"4a",x"a3"),
   936 => (x"12",x"4a",x"a3",x"d4"),
   937 => (x"4a",x"a3",x"d6",x"51"),
   938 => (x"a3",x"d8",x"51",x"12"),
   939 => (x"dc",x"51",x"12",x"4a"),
   940 => (x"51",x"12",x"4a",x"a3"),
   941 => (x"12",x"4a",x"a3",x"de"),
   942 => (x"c0",x"7e",x"c1",x"51"),
   943 => (x"49",x"74",x"87",x"fc"),
   944 => (x"c0",x"05",x"99",x"c8"),
   945 => (x"49",x"74",x"87",x"ed"),
   946 => (x"d3",x"05",x"99",x"d0"),
   947 => (x"66",x"e0",x"c0",x"87"),
   948 => (x"87",x"cc",x"c0",x"02"),
   949 => (x"e0",x"c0",x"49",x"73"),
   950 => (x"98",x"70",x"0f",x"66"),
   951 => (x"87",x"d3",x"c0",x"02"),
   952 => (x"c6",x"c0",x"05",x"6e"),
   953 => (x"e4",x"f2",x"c2",x"87"),
   954 => (x"c0",x"50",x"c0",x"48"),
   955 => (x"48",x"bf",x"ec",x"fe"),
   956 => (x"c2",x"87",x"e9",x"c2"),
   957 => (x"c0",x"48",x"f1",x"f2"),
   958 => (x"f2",x"c2",x"7e",x"50"),
   959 => (x"c2",x"49",x"bf",x"e0"),
   960 => (x"4a",x"bf",x"d0",x"ea"),
   961 => (x"fb",x"04",x"aa",x"71"),
   962 => (x"ff",x"cf",x"87",x"f4"),
   963 => (x"4c",x"f8",x"ff",x"ff"),
   964 => (x"bf",x"c4",x"f7",x"c2"),
   965 => (x"87",x"c8",x"c0",x"05"),
   966 => (x"bf",x"dc",x"f2",x"c2"),
   967 => (x"87",x"fa",x"c1",x"02"),
   968 => (x"bf",x"cc",x"ea",x"c2"),
   969 => (x"87",x"fa",x"e6",x"49"),
   970 => (x"58",x"d0",x"ea",x"c2"),
   971 => (x"c2",x"48",x"a6",x"c4"),
   972 => (x"78",x"bf",x"cc",x"ea"),
   973 => (x"bf",x"dc",x"f2",x"c2"),
   974 => (x"87",x"db",x"c0",x"02"),
   975 => (x"74",x"49",x"66",x"c4"),
   976 => (x"02",x"a9",x"74",x"99"),
   977 => (x"c8",x"87",x"c8",x"c0"),
   978 => (x"78",x"c0",x"48",x"a6"),
   979 => (x"c8",x"87",x"e7",x"c0"),
   980 => (x"78",x"c1",x"48",x"a6"),
   981 => (x"c4",x"87",x"df",x"c0"),
   982 => (x"ff",x"cf",x"49",x"66"),
   983 => (x"02",x"a9",x"99",x"f8"),
   984 => (x"cc",x"87",x"c8",x"c0"),
   985 => (x"78",x"c0",x"48",x"a6"),
   986 => (x"cc",x"87",x"c5",x"c0"),
   987 => (x"78",x"c1",x"48",x"a6"),
   988 => (x"cc",x"48",x"a6",x"c8"),
   989 => (x"66",x"c8",x"78",x"66"),
   990 => (x"87",x"de",x"c0",x"05"),
   991 => (x"c2",x"49",x"66",x"c4"),
   992 => (x"d4",x"f2",x"c2",x"89"),
   993 => (x"f6",x"c2",x"91",x"bf"),
   994 => (x"71",x"48",x"bf",x"f0"),
   995 => (x"cc",x"ea",x"c2",x"80"),
   996 => (x"d0",x"ea",x"c2",x"58"),
   997 => (x"f9",x"78",x"c0",x"48"),
   998 => (x"48",x"c0",x"87",x"d4"),
   999 => (x"ff",x"ff",x"ff",x"cf"),
  1000 => (x"8e",x"f0",x"4c",x"f8"),
  1001 => (x"4c",x"26",x"4d",x"26"),
  1002 => (x"4f",x"26",x"4b",x"26"),
  1003 => (x"00",x"00",x"00",x"00"),
  1004 => (x"ff",x"ff",x"ff",x"ff"),
  1005 => (x"00",x"00",x"0f",x"bc"),
  1006 => (x"00",x"00",x"0f",x"c8"),
  1007 => (x"33",x"54",x"41",x"46"),
  1008 => (x"20",x"20",x"20",x"32"),
  1009 => (x"00",x"00",x"00",x"00"),
  1010 => (x"31",x"54",x"41",x"46"),
  1011 => (x"20",x"20",x"20",x"36"),
  1012 => (x"d4",x"ff",x"1e",x"00"),
  1013 => (x"78",x"ff",x"c3",x"48"),
  1014 => (x"4f",x"26",x"48",x"68"),
  1015 => (x"48",x"d4",x"ff",x"1e"),
  1016 => (x"ff",x"78",x"ff",x"c3"),
  1017 => (x"e1",x"c0",x"48",x"d0"),
  1018 => (x"48",x"d4",x"ff",x"78"),
  1019 => (x"4f",x"26",x"78",x"d4"),
  1020 => (x"48",x"d0",x"ff",x"1e"),
  1021 => (x"26",x"78",x"e0",x"c0"),
  1022 => (x"d4",x"ff",x"1e",x"4f"),
  1023 => (x"99",x"49",x"70",x"87"),
  1024 => (x"c0",x"87",x"c6",x"02"),
  1025 => (x"f1",x"05",x"a9",x"fb"),
  1026 => (x"26",x"48",x"71",x"87"),
  1027 => (x"5b",x"5e",x"0e",x"4f"),
  1028 => (x"4b",x"71",x"0e",x"5c"),
  1029 => (x"f8",x"fe",x"4c",x"c0"),
  1030 => (x"99",x"49",x"70",x"87"),
  1031 => (x"87",x"f9",x"c0",x"02"),
  1032 => (x"02",x"a9",x"ec",x"c0"),
  1033 => (x"c0",x"87",x"f2",x"c0"),
  1034 => (x"c0",x"02",x"a9",x"fb"),
  1035 => (x"66",x"cc",x"87",x"eb"),
  1036 => (x"c7",x"03",x"ac",x"b7"),
  1037 => (x"02",x"66",x"d0",x"87"),
  1038 => (x"53",x"71",x"87",x"c2"),
  1039 => (x"c2",x"02",x"99",x"71"),
  1040 => (x"fe",x"84",x"c1",x"87"),
  1041 => (x"49",x"70",x"87",x"cb"),
  1042 => (x"87",x"cd",x"02",x"99"),
  1043 => (x"02",x"a9",x"ec",x"c0"),
  1044 => (x"fb",x"c0",x"87",x"c7"),
  1045 => (x"d5",x"ff",x"05",x"a9"),
  1046 => (x"02",x"66",x"d0",x"87"),
  1047 => (x"97",x"c0",x"87",x"c3"),
  1048 => (x"a9",x"ec",x"c0",x"7b"),
  1049 => (x"74",x"87",x"c4",x"05"),
  1050 => (x"74",x"87",x"c5",x"4a"),
  1051 => (x"8a",x"0a",x"c0",x"4a"),
  1052 => (x"4c",x"26",x"48",x"72"),
  1053 => (x"4f",x"26",x"4b",x"26"),
  1054 => (x"87",x"d5",x"fd",x"1e"),
  1055 => (x"f0",x"c0",x"49",x"70"),
  1056 => (x"87",x"c9",x"04",x"a9"),
  1057 => (x"01",x"a9",x"f9",x"c0"),
  1058 => (x"f0",x"c0",x"87",x"c3"),
  1059 => (x"a9",x"c1",x"c1",x"89"),
  1060 => (x"c1",x"87",x"c9",x"04"),
  1061 => (x"c3",x"01",x"a9",x"da"),
  1062 => (x"89",x"f7",x"c0",x"87"),
  1063 => (x"4f",x"26",x"48",x"71"),
  1064 => (x"5c",x"5b",x"5e",x"0e"),
  1065 => (x"86",x"f8",x"0e",x"5d"),
  1066 => (x"7e",x"c0",x"4c",x"71"),
  1067 => (x"c0",x"87",x"ed",x"fc"),
  1068 => (x"c0",x"c5",x"c1",x"4b"),
  1069 => (x"c0",x"49",x"bf",x"97"),
  1070 => (x"87",x"cf",x"04",x"a9"),
  1071 => (x"c1",x"87",x"fa",x"fc"),
  1072 => (x"c0",x"c5",x"c1",x"83"),
  1073 => (x"ab",x"49",x"bf",x"97"),
  1074 => (x"c1",x"87",x"f1",x"06"),
  1075 => (x"bf",x"97",x"c0",x"c5"),
  1076 => (x"fb",x"87",x"cf",x"02"),
  1077 => (x"49",x"70",x"87",x"fb"),
  1078 => (x"87",x"c6",x"02",x"99"),
  1079 => (x"05",x"a9",x"ec",x"c0"),
  1080 => (x"4b",x"c0",x"87",x"f1"),
  1081 => (x"70",x"87",x"ea",x"fb"),
  1082 => (x"87",x"e5",x"fb",x"4d"),
  1083 => (x"fb",x"58",x"a6",x"c8"),
  1084 => (x"4a",x"70",x"87",x"df"),
  1085 => (x"a4",x"c8",x"83",x"c1"),
  1086 => (x"49",x"69",x"97",x"49"),
  1087 => (x"87",x"da",x"05",x"ad"),
  1088 => (x"97",x"49",x"a4",x"c9"),
  1089 => (x"66",x"c4",x"49",x"69"),
  1090 => (x"87",x"ce",x"05",x"a9"),
  1091 => (x"97",x"49",x"a4",x"ca"),
  1092 => (x"05",x"aa",x"49",x"69"),
  1093 => (x"7e",x"c1",x"87",x"c4"),
  1094 => (x"ec",x"c0",x"87",x"d0"),
  1095 => (x"87",x"c6",x"02",x"ad"),
  1096 => (x"05",x"ad",x"fb",x"c0"),
  1097 => (x"4b",x"c0",x"87",x"c4"),
  1098 => (x"02",x"6e",x"7e",x"c1"),
  1099 => (x"fa",x"87",x"f5",x"fe"),
  1100 => (x"48",x"73",x"87",x"fe"),
  1101 => (x"4d",x"26",x"8e",x"f8"),
  1102 => (x"4b",x"26",x"4c",x"26"),
  1103 => (x"00",x"00",x"4f",x"26"),
  1104 => (x"1e",x"73",x"1e",x"00"),
  1105 => (x"c8",x"4b",x"d4",x"ff"),
  1106 => (x"d0",x"ff",x"4a",x"66"),
  1107 => (x"78",x"c5",x"c8",x"48"),
  1108 => (x"c1",x"48",x"d4",x"ff"),
  1109 => (x"7b",x"11",x"78",x"d4"),
  1110 => (x"f9",x"05",x"8a",x"c1"),
  1111 => (x"48",x"d0",x"ff",x"87"),
  1112 => (x"4b",x"26",x"78",x"c4"),
  1113 => (x"5e",x"0e",x"4f",x"26"),
  1114 => (x"0e",x"5d",x"5c",x"5b"),
  1115 => (x"7e",x"71",x"86",x"f8"),
  1116 => (x"f7",x"c2",x"1e",x"6e"),
  1117 => (x"df",x"ff",x"49",x"d4"),
  1118 => (x"86",x"c4",x"87",x"df"),
  1119 => (x"c4",x"02",x"98",x"70"),
  1120 => (x"f4",x"c1",x"87",x"e4"),
  1121 => (x"6e",x"4c",x"bf",x"c8"),
  1122 => (x"87",x"d4",x"fc",x"49"),
  1123 => (x"70",x"58",x"a6",x"c8"),
  1124 => (x"87",x"c5",x"05",x"98"),
  1125 => (x"c1",x"48",x"a6",x"c4"),
  1126 => (x"48",x"d0",x"ff",x"78"),
  1127 => (x"d4",x"ff",x"78",x"c5"),
  1128 => (x"78",x"d5",x"c1",x"48"),
  1129 => (x"c1",x"49",x"66",x"c4"),
  1130 => (x"c1",x"31",x"c6",x"89"),
  1131 => (x"bf",x"97",x"c0",x"f4"),
  1132 => (x"b0",x"71",x"48",x"4a"),
  1133 => (x"78",x"08",x"d4",x"ff"),
  1134 => (x"c4",x"48",x"d0",x"ff"),
  1135 => (x"d0",x"f7",x"c2",x"78"),
  1136 => (x"d0",x"49",x"bf",x"97"),
  1137 => (x"87",x"dd",x"02",x"99"),
  1138 => (x"d4",x"ff",x"78",x"c5"),
  1139 => (x"78",x"d6",x"c1",x"48"),
  1140 => (x"d4",x"ff",x"4a",x"c0"),
  1141 => (x"78",x"ff",x"c3",x"48"),
  1142 => (x"e0",x"c0",x"82",x"c1"),
  1143 => (x"87",x"f2",x"04",x"aa"),
  1144 => (x"c4",x"48",x"d0",x"ff"),
  1145 => (x"48",x"d4",x"ff",x"78"),
  1146 => (x"ff",x"78",x"ff",x"c3"),
  1147 => (x"78",x"c5",x"48",x"d0"),
  1148 => (x"c1",x"48",x"d4",x"ff"),
  1149 => (x"78",x"c1",x"78",x"d3"),
  1150 => (x"c4",x"48",x"d0",x"ff"),
  1151 => (x"ac",x"b7",x"c0",x"78"),
  1152 => (x"87",x"cb",x"c2",x"06"),
  1153 => (x"bf",x"dc",x"f7",x"c2"),
  1154 => (x"7e",x"74",x"8c",x"4b"),
  1155 => (x"c1",x"02",x"9b",x"73"),
  1156 => (x"c0",x"c8",x"87",x"dd"),
  1157 => (x"b7",x"c0",x"8b",x"4d"),
  1158 => (x"87",x"c6",x"03",x"ab"),
  1159 => (x"4d",x"a3",x"c0",x"c8"),
  1160 => (x"f7",x"c2",x"4b",x"c0"),
  1161 => (x"49",x"bf",x"97",x"d0"),
  1162 => (x"cf",x"02",x"99",x"d0"),
  1163 => (x"c2",x"1e",x"c0",x"87"),
  1164 => (x"e2",x"49",x"d4",x"f7"),
  1165 => (x"86",x"c4",x"87",x"e1"),
  1166 => (x"87",x"d8",x"4c",x"70"),
  1167 => (x"1e",x"d4",x"ea",x"c2"),
  1168 => (x"49",x"d4",x"f7",x"c2"),
  1169 => (x"70",x"87",x"d0",x"e2"),
  1170 => (x"c2",x"1e",x"75",x"4c"),
  1171 => (x"fb",x"49",x"d4",x"ea"),
  1172 => (x"86",x"c8",x"87",x"ef"),
  1173 => (x"c5",x"05",x"9c",x"74"),
  1174 => (x"c1",x"48",x"c0",x"87"),
  1175 => (x"1e",x"c1",x"87",x"ca"),
  1176 => (x"49",x"d4",x"f7",x"c2"),
  1177 => (x"c4",x"87",x"d5",x"e0"),
  1178 => (x"05",x"9b",x"73",x"86"),
  1179 => (x"6e",x"87",x"e3",x"fe"),
  1180 => (x"ac",x"b7",x"c0",x"4c"),
  1181 => (x"c2",x"87",x"d1",x"06"),
  1182 => (x"c0",x"48",x"d4",x"f7"),
  1183 => (x"c0",x"80",x"d0",x"78"),
  1184 => (x"c2",x"80",x"f4",x"78"),
  1185 => (x"78",x"bf",x"e0",x"f7"),
  1186 => (x"01",x"ac",x"b7",x"c0"),
  1187 => (x"ff",x"87",x"f5",x"fd"),
  1188 => (x"78",x"c5",x"48",x"d0"),
  1189 => (x"c1",x"48",x"d4",x"ff"),
  1190 => (x"78",x"c0",x"78",x"d3"),
  1191 => (x"c4",x"48",x"d0",x"ff"),
  1192 => (x"c0",x"48",x"c1",x"78"),
  1193 => (x"48",x"c0",x"87",x"c2"),
  1194 => (x"4d",x"26",x"8e",x"f8"),
  1195 => (x"4b",x"26",x"4c",x"26"),
  1196 => (x"5e",x"0e",x"4f",x"26"),
  1197 => (x"0e",x"5d",x"5c",x"5b"),
  1198 => (x"4d",x"71",x"86",x"fc"),
  1199 => (x"ad",x"4c",x"4b",x"c0"),
  1200 => (x"87",x"e8",x"c0",x"04"),
  1201 => (x"1e",x"e0",x"c2",x"c1"),
  1202 => (x"c4",x"02",x"9c",x"74"),
  1203 => (x"c2",x"4a",x"c0",x"87"),
  1204 => (x"72",x"4a",x"c1",x"87"),
  1205 => (x"87",x"e0",x"eb",x"49"),
  1206 => (x"7e",x"70",x"86",x"c4"),
  1207 => (x"05",x"6e",x"83",x"c1"),
  1208 => (x"4b",x"75",x"87",x"c2"),
  1209 => (x"ab",x"75",x"84",x"c1"),
  1210 => (x"87",x"d8",x"ff",x"06"),
  1211 => (x"8e",x"fc",x"48",x"6e"),
  1212 => (x"4c",x"26",x"4d",x"26"),
  1213 => (x"4f",x"26",x"4b",x"26"),
  1214 => (x"5c",x"5b",x"5e",x"0e"),
  1215 => (x"cc",x"4b",x"71",x"0e"),
  1216 => (x"87",x"d8",x"02",x"66"),
  1217 => (x"8c",x"f0",x"c0",x"4c"),
  1218 => (x"74",x"87",x"d8",x"02"),
  1219 => (x"02",x"8a",x"c1",x"4a"),
  1220 => (x"02",x"8a",x"87",x"d1"),
  1221 => (x"02",x"8a",x"87",x"cd"),
  1222 => (x"87",x"d9",x"87",x"c9"),
  1223 => (x"c5",x"f9",x"49",x"73"),
  1224 => (x"74",x"87",x"d2",x"87"),
  1225 => (x"c1",x"49",x"c0",x"1e"),
  1226 => (x"74",x"87",x"fd",x"d9"),
  1227 => (x"c1",x"49",x"73",x"1e"),
  1228 => (x"c8",x"87",x"f5",x"d9"),
  1229 => (x"26",x"4c",x"26",x"86"),
  1230 => (x"0e",x"4f",x"26",x"4b"),
  1231 => (x"5d",x"5c",x"5b",x"5e"),
  1232 => (x"71",x"86",x"fc",x"0e"),
  1233 => (x"91",x"de",x"49",x"4c"),
  1234 => (x"4d",x"f4",x"f8",x"c2"),
  1235 => (x"6d",x"97",x"85",x"71"),
  1236 => (x"87",x"dc",x"c1",x"02"),
  1237 => (x"bf",x"e4",x"f8",x"c2"),
  1238 => (x"71",x"81",x"74",x"49"),
  1239 => (x"70",x"87",x"d3",x"fd"),
  1240 => (x"02",x"98",x"48",x"7e"),
  1241 => (x"c2",x"87",x"f2",x"c0"),
  1242 => (x"70",x"4b",x"e8",x"f8"),
  1243 => (x"fe",x"49",x"cb",x"4a"),
  1244 => (x"74",x"87",x"f1",x"f6"),
  1245 => (x"c1",x"93",x"cc",x"4b"),
  1246 => (x"c4",x"83",x"cc",x"f4"),
  1247 => (x"fc",x"ce",x"c1",x"83"),
  1248 => (x"c1",x"49",x"74",x"7b"),
  1249 => (x"75",x"87",x"e9",x"c4"),
  1250 => (x"c4",x"f4",x"c1",x"7b"),
  1251 => (x"1e",x"49",x"bf",x"97"),
  1252 => (x"49",x"e8",x"f8",x"c2"),
  1253 => (x"c4",x"87",x"e1",x"fd"),
  1254 => (x"c1",x"49",x"74",x"86"),
  1255 => (x"c0",x"87",x"d1",x"c4"),
  1256 => (x"ec",x"c5",x"c1",x"49"),
  1257 => (x"cc",x"f7",x"c2",x"87"),
  1258 => (x"49",x"50",x"c0",x"48"),
  1259 => (x"87",x"cb",x"e2",x"c0"),
  1260 => (x"4d",x"26",x"8e",x"fc"),
  1261 => (x"4b",x"26",x"4c",x"26"),
  1262 => (x"00",x"00",x"4f",x"26"),
  1263 => (x"64",x"61",x"6f",x"4c"),
  1264 => (x"2e",x"67",x"6e",x"69"),
  1265 => (x"1e",x"00",x"2e",x"2e"),
  1266 => (x"4b",x"71",x"1e",x"73"),
  1267 => (x"e4",x"f8",x"c2",x"49"),
  1268 => (x"fb",x"71",x"81",x"bf"),
  1269 => (x"4a",x"70",x"87",x"dc"),
  1270 => (x"87",x"c4",x"02",x"9a"),
  1271 => (x"87",x"de",x"e6",x"49"),
  1272 => (x"48",x"e4",x"f8",x"c2"),
  1273 => (x"49",x"73",x"78",x"c0"),
  1274 => (x"26",x"87",x"fa",x"c1"),
  1275 => (x"1e",x"4f",x"26",x"4b"),
  1276 => (x"4b",x"71",x"1e",x"73"),
  1277 => (x"02",x"4a",x"a3",x"c4"),
  1278 => (x"c1",x"87",x"d0",x"c1"),
  1279 => (x"87",x"dc",x"02",x"8a"),
  1280 => (x"f2",x"c0",x"02",x"8a"),
  1281 => (x"c1",x"05",x"8a",x"87"),
  1282 => (x"f8",x"c2",x"87",x"d3"),
  1283 => (x"c1",x"02",x"bf",x"e4"),
  1284 => (x"c1",x"48",x"87",x"cb"),
  1285 => (x"e8",x"f8",x"c2",x"88"),
  1286 => (x"87",x"c1",x"c1",x"58"),
  1287 => (x"bf",x"e4",x"f8",x"c2"),
  1288 => (x"c2",x"89",x"c6",x"49"),
  1289 => (x"c0",x"59",x"e8",x"f8"),
  1290 => (x"c0",x"03",x"a9",x"b7"),
  1291 => (x"f8",x"c2",x"87",x"ef"),
  1292 => (x"78",x"c0",x"48",x"e4"),
  1293 => (x"c2",x"87",x"e6",x"c0"),
  1294 => (x"02",x"bf",x"e0",x"f8"),
  1295 => (x"f8",x"c2",x"87",x"df"),
  1296 => (x"c1",x"48",x"bf",x"e4"),
  1297 => (x"e8",x"f8",x"c2",x"80"),
  1298 => (x"c2",x"87",x"d2",x"58"),
  1299 => (x"02",x"bf",x"e0",x"f8"),
  1300 => (x"f8",x"c2",x"87",x"cb"),
  1301 => (x"c6",x"48",x"bf",x"e4"),
  1302 => (x"e8",x"f8",x"c2",x"80"),
  1303 => (x"c4",x"49",x"73",x"58"),
  1304 => (x"26",x"4b",x"26",x"87"),
  1305 => (x"5b",x"5e",x"0e",x"4f"),
  1306 => (x"f0",x"0e",x"5d",x"5c"),
  1307 => (x"59",x"a6",x"d0",x"86"),
  1308 => (x"4d",x"d4",x"ea",x"c2"),
  1309 => (x"f8",x"c2",x"4c",x"c0"),
  1310 => (x"78",x"c1",x"48",x"e0"),
  1311 => (x"c0",x"48",x"a6",x"c8"),
  1312 => (x"c2",x"7e",x"75",x"78"),
  1313 => (x"48",x"bf",x"e4",x"f8"),
  1314 => (x"c1",x"06",x"a8",x"c0"),
  1315 => (x"a6",x"c8",x"87",x"c0"),
  1316 => (x"c2",x"7e",x"75",x"5c"),
  1317 => (x"98",x"48",x"d4",x"ea"),
  1318 => (x"87",x"f2",x"c0",x"02"),
  1319 => (x"c1",x"4d",x"66",x"c4"),
  1320 => (x"cc",x"1e",x"e0",x"c2"),
  1321 => (x"87",x"c4",x"02",x"66"),
  1322 => (x"87",x"c2",x"4c",x"c0"),
  1323 => (x"49",x"74",x"4c",x"c1"),
  1324 => (x"c4",x"87",x"c5",x"e4"),
  1325 => (x"c1",x"7e",x"70",x"86"),
  1326 => (x"48",x"66",x"c8",x"85"),
  1327 => (x"a6",x"cc",x"80",x"c1"),
  1328 => (x"e4",x"f8",x"c2",x"58"),
  1329 => (x"c5",x"03",x"ad",x"bf"),
  1330 => (x"ff",x"05",x"6e",x"87"),
  1331 => (x"4d",x"6e",x"87",x"d1"),
  1332 => (x"9d",x"75",x"4c",x"c0"),
  1333 => (x"87",x"dc",x"c3",x"02"),
  1334 => (x"1e",x"e0",x"c2",x"c1"),
  1335 => (x"c7",x"02",x"66",x"cc"),
  1336 => (x"48",x"a6",x"c8",x"87"),
  1337 => (x"87",x"c5",x"78",x"c0"),
  1338 => (x"c1",x"48",x"a6",x"c8"),
  1339 => (x"49",x"66",x"c8",x"78"),
  1340 => (x"c4",x"87",x"c5",x"e3"),
  1341 => (x"48",x"7e",x"70",x"86"),
  1342 => (x"e4",x"c2",x"02",x"98"),
  1343 => (x"81",x"cb",x"49",x"87"),
  1344 => (x"d0",x"49",x"69",x"97"),
  1345 => (x"d4",x"c1",x"02",x"99"),
  1346 => (x"cc",x"49",x"74",x"87"),
  1347 => (x"cc",x"f4",x"c1",x"91"),
  1348 => (x"c7",x"cf",x"c1",x"81"),
  1349 => (x"c3",x"81",x"c8",x"79"),
  1350 => (x"49",x"74",x"51",x"ff"),
  1351 => (x"f8",x"c2",x"91",x"de"),
  1352 => (x"85",x"71",x"4d",x"f4"),
  1353 => (x"7d",x"97",x"c1",x"c2"),
  1354 => (x"c0",x"49",x"a5",x"c1"),
  1355 => (x"f2",x"c2",x"51",x"e0"),
  1356 => (x"02",x"bf",x"97",x"e4"),
  1357 => (x"84",x"c1",x"87",x"d2"),
  1358 => (x"c2",x"4b",x"a5",x"c2"),
  1359 => (x"db",x"4a",x"e4",x"f2"),
  1360 => (x"df",x"ef",x"fe",x"49"),
  1361 => (x"87",x"d9",x"c1",x"87"),
  1362 => (x"c0",x"49",x"a5",x"cd"),
  1363 => (x"c2",x"84",x"c1",x"51"),
  1364 => (x"4a",x"6e",x"4b",x"a5"),
  1365 => (x"ef",x"fe",x"49",x"cb"),
  1366 => (x"c4",x"c1",x"87",x"ca"),
  1367 => (x"cc",x"49",x"74",x"87"),
  1368 => (x"cc",x"f4",x"c1",x"91"),
  1369 => (x"fb",x"cc",x"c1",x"81"),
  1370 => (x"e4",x"f2",x"c2",x"79"),
  1371 => (x"d8",x"02",x"bf",x"97"),
  1372 => (x"de",x"49",x"74",x"87"),
  1373 => (x"c2",x"84",x"c1",x"91"),
  1374 => (x"71",x"4b",x"f4",x"f8"),
  1375 => (x"e4",x"f2",x"c2",x"83"),
  1376 => (x"fe",x"49",x"dd",x"4a"),
  1377 => (x"d8",x"87",x"dd",x"ee"),
  1378 => (x"de",x"4b",x"74",x"87"),
  1379 => (x"f4",x"f8",x"c2",x"93"),
  1380 => (x"49",x"a3",x"cb",x"83"),
  1381 => (x"84",x"c1",x"51",x"c0"),
  1382 => (x"cb",x"4a",x"6e",x"73"),
  1383 => (x"c3",x"ee",x"fe",x"49"),
  1384 => (x"48",x"66",x"c8",x"87"),
  1385 => (x"a6",x"cc",x"80",x"c1"),
  1386 => (x"03",x"ac",x"c7",x"58"),
  1387 => (x"6e",x"87",x"c5",x"c0"),
  1388 => (x"87",x"e4",x"fc",x"05"),
  1389 => (x"c0",x"03",x"ac",x"c7"),
  1390 => (x"f8",x"c2",x"87",x"e4"),
  1391 => (x"78",x"c0",x"48",x"e0"),
  1392 => (x"91",x"cc",x"49",x"74"),
  1393 => (x"81",x"cc",x"f4",x"c1"),
  1394 => (x"79",x"fb",x"cc",x"c1"),
  1395 => (x"91",x"de",x"49",x"74"),
  1396 => (x"81",x"f4",x"f8",x"c2"),
  1397 => (x"84",x"c1",x"51",x"c0"),
  1398 => (x"ff",x"04",x"ac",x"c7"),
  1399 => (x"f5",x"c1",x"87",x"dc"),
  1400 => (x"50",x"c0",x"48",x"e8"),
  1401 => (x"d9",x"c1",x"80",x"f7"),
  1402 => (x"d8",x"c1",x"40",x"d5"),
  1403 => (x"80",x"c8",x"78",x"c8"),
  1404 => (x"78",x"ef",x"cf",x"c1"),
  1405 => (x"c0",x"49",x"66",x"cc"),
  1406 => (x"f0",x"87",x"f5",x"fa"),
  1407 => (x"26",x"4d",x"26",x"8e"),
  1408 => (x"26",x"4b",x"26",x"4c"),
  1409 => (x"00",x"00",x"00",x"4f"),
  1410 => (x"61",x"42",x"20",x"80"),
  1411 => (x"1e",x"00",x"6b",x"63"),
  1412 => (x"4b",x"71",x"1e",x"73"),
  1413 => (x"c1",x"91",x"cc",x"49"),
  1414 => (x"c8",x"81",x"cc",x"f4"),
  1415 => (x"f4",x"c1",x"4a",x"a1"),
  1416 => (x"50",x"12",x"48",x"c0"),
  1417 => (x"c1",x"4a",x"a1",x"c9"),
  1418 => (x"12",x"48",x"c0",x"c5"),
  1419 => (x"c1",x"81",x"ca",x"50"),
  1420 => (x"11",x"48",x"c4",x"f4"),
  1421 => (x"c4",x"f4",x"c1",x"50"),
  1422 => (x"1e",x"49",x"bf",x"97"),
  1423 => (x"f7",x"f2",x"49",x"c0"),
  1424 => (x"f8",x"49",x"73",x"87"),
  1425 => (x"8e",x"fc",x"87",x"df"),
  1426 => (x"4f",x"26",x"4b",x"26"),
  1427 => (x"c0",x"49",x"c0",x"1e"),
  1428 => (x"26",x"87",x"fe",x"fa"),
  1429 => (x"4a",x"71",x"1e",x"4f"),
  1430 => (x"c1",x"91",x"cc",x"49"),
  1431 => (x"c8",x"81",x"cc",x"f4"),
  1432 => (x"cc",x"f7",x"c2",x"81"),
  1433 => (x"c0",x"50",x"11",x"48"),
  1434 => (x"fe",x"49",x"a2",x"f0"),
  1435 => (x"c0",x"87",x"dd",x"e8"),
  1436 => (x"87",x"c7",x"d7",x"49"),
  1437 => (x"ff",x"1e",x"4f",x"26"),
  1438 => (x"ff",x"c3",x"4a",x"d4"),
  1439 => (x"48",x"d0",x"ff",x"7a"),
  1440 => (x"de",x"78",x"e1",x"c0"),
  1441 => (x"48",x"7a",x"71",x"7a"),
  1442 => (x"70",x"28",x"b7",x"c8"),
  1443 => (x"d0",x"48",x"71",x"7a"),
  1444 => (x"7a",x"70",x"28",x"b7"),
  1445 => (x"b7",x"d8",x"48",x"71"),
  1446 => (x"ff",x"7a",x"70",x"28"),
  1447 => (x"e0",x"c0",x"48",x"d0"),
  1448 => (x"0e",x"4f",x"26",x"78"),
  1449 => (x"5d",x"5c",x"5b",x"5e"),
  1450 => (x"71",x"86",x"f4",x"0e"),
  1451 => (x"91",x"cc",x"49",x"4d"),
  1452 => (x"81",x"cc",x"f4",x"c1"),
  1453 => (x"ca",x"4a",x"a1",x"c8"),
  1454 => (x"a6",x"c4",x"7e",x"a1"),
  1455 => (x"c8",x"f7",x"c2",x"48"),
  1456 => (x"97",x"6e",x"78",x"bf"),
  1457 => (x"66",x"c4",x"4b",x"bf"),
  1458 => (x"12",x"2c",x"73",x"4c"),
  1459 => (x"58",x"a6",x"cc",x"48"),
  1460 => (x"84",x"c1",x"9c",x"70"),
  1461 => (x"69",x"97",x"81",x"c9"),
  1462 => (x"04",x"ac",x"b7",x"49"),
  1463 => (x"4c",x"c0",x"87",x"c2"),
  1464 => (x"4a",x"bf",x"97",x"6e"),
  1465 => (x"72",x"49",x"66",x"c8"),
  1466 => (x"c4",x"b9",x"ff",x"31"),
  1467 => (x"48",x"74",x"99",x"66"),
  1468 => (x"4a",x"70",x"30",x"72"),
  1469 => (x"cc",x"f7",x"c2",x"b1"),
  1470 => (x"f9",x"fd",x"71",x"59"),
  1471 => (x"c2",x"1e",x"c7",x"87"),
  1472 => (x"1e",x"bf",x"dc",x"f8"),
  1473 => (x"1e",x"cc",x"f4",x"c1"),
  1474 => (x"97",x"cc",x"f7",x"c2"),
  1475 => (x"f4",x"c1",x"49",x"bf"),
  1476 => (x"c0",x"49",x"75",x"87"),
  1477 => (x"e8",x"87",x"d9",x"f6"),
  1478 => (x"26",x"4d",x"26",x"8e"),
  1479 => (x"26",x"4b",x"26",x"4c"),
  1480 => (x"1e",x"73",x"1e",x"4f"),
  1481 => (x"fd",x"49",x"4b",x"71"),
  1482 => (x"49",x"73",x"87",x"f9"),
  1483 => (x"26",x"87",x"f4",x"fd"),
  1484 => (x"1e",x"4f",x"26",x"4b"),
  1485 => (x"4b",x"71",x"1e",x"73"),
  1486 => (x"02",x"4a",x"a3",x"c2"),
  1487 => (x"8a",x"c1",x"87",x"d6"),
  1488 => (x"87",x"e2",x"c0",x"05"),
  1489 => (x"bf",x"dc",x"f8",x"c2"),
  1490 => (x"48",x"87",x"db",x"02"),
  1491 => (x"f8",x"c2",x"88",x"c1"),
  1492 => (x"87",x"d2",x"58",x"e0"),
  1493 => (x"bf",x"e0",x"f8",x"c2"),
  1494 => (x"c2",x"87",x"cb",x"02"),
  1495 => (x"48",x"bf",x"dc",x"f8"),
  1496 => (x"f8",x"c2",x"80",x"c1"),
  1497 => (x"1e",x"c7",x"58",x"e0"),
  1498 => (x"bf",x"dc",x"f8",x"c2"),
  1499 => (x"cc",x"f4",x"c1",x"1e"),
  1500 => (x"cc",x"f7",x"c2",x"1e"),
  1501 => (x"cc",x"49",x"bf",x"97"),
  1502 => (x"c0",x"49",x"73",x"87"),
  1503 => (x"f4",x"87",x"f1",x"f4"),
  1504 => (x"26",x"4b",x"26",x"8e"),
  1505 => (x"5b",x"5e",x"0e",x"4f"),
  1506 => (x"ff",x"0e",x"5d",x"5c"),
  1507 => (x"e4",x"c0",x"86",x"cc"),
  1508 => (x"a6",x"cc",x"59",x"a6"),
  1509 => (x"c4",x"78",x"c0",x"48"),
  1510 => (x"c4",x"78",x"c0",x"80"),
  1511 => (x"66",x"c8",x"c1",x"80"),
  1512 => (x"c1",x"80",x"c4",x"78"),
  1513 => (x"c1",x"80",x"c4",x"78"),
  1514 => (x"e0",x"f8",x"c2",x"78"),
  1515 => (x"e0",x"78",x"c1",x"48"),
  1516 => (x"c4",x"e1",x"87",x"ea"),
  1517 => (x"87",x"d9",x"e0",x"87"),
  1518 => (x"fb",x"c0",x"4c",x"70"),
  1519 => (x"f3",x"c1",x"02",x"ac"),
  1520 => (x"66",x"e0",x"c0",x"87"),
  1521 => (x"87",x"e8",x"c1",x"05"),
  1522 => (x"4a",x"66",x"c4",x"c1"),
  1523 => (x"7e",x"6a",x"82",x"c4"),
  1524 => (x"48",x"dc",x"f0",x"c1"),
  1525 => (x"41",x"20",x"49",x"6e"),
  1526 => (x"51",x"10",x"41",x"20"),
  1527 => (x"48",x"66",x"c4",x"c1"),
  1528 => (x"78",x"cf",x"d8",x"c1"),
  1529 => (x"81",x"c7",x"49",x"6a"),
  1530 => (x"c4",x"c1",x"51",x"74"),
  1531 => (x"81",x"c8",x"49",x"66"),
  1532 => (x"a6",x"d8",x"51",x"c1"),
  1533 => (x"c1",x"78",x"c2",x"48"),
  1534 => (x"c9",x"49",x"66",x"c4"),
  1535 => (x"c1",x"51",x"c0",x"81"),
  1536 => (x"ca",x"49",x"66",x"c4"),
  1537 => (x"c1",x"51",x"c0",x"81"),
  1538 => (x"6a",x"1e",x"d8",x"1e"),
  1539 => (x"ff",x"81",x"c8",x"49"),
  1540 => (x"c8",x"87",x"fa",x"df"),
  1541 => (x"66",x"c8",x"c1",x"86"),
  1542 => (x"01",x"a8",x"c0",x"48"),
  1543 => (x"a6",x"d0",x"87",x"c7"),
  1544 => (x"cf",x"78",x"c1",x"48"),
  1545 => (x"66",x"c8",x"c1",x"87"),
  1546 => (x"d8",x"88",x"c1",x"48"),
  1547 => (x"87",x"c4",x"58",x"a6"),
  1548 => (x"87",x"c5",x"df",x"ff"),
  1549 => (x"cd",x"02",x"9c",x"74"),
  1550 => (x"66",x"d0",x"87",x"d9"),
  1551 => (x"66",x"cc",x"c1",x"48"),
  1552 => (x"ce",x"cd",x"03",x"a8"),
  1553 => (x"48",x"a6",x"c8",x"87"),
  1554 => (x"ff",x"7e",x"78",x"c0"),
  1555 => (x"70",x"87",x"c2",x"de"),
  1556 => (x"ac",x"d0",x"c1",x"4c"),
  1557 => (x"87",x"e7",x"c2",x"05"),
  1558 => (x"6e",x"48",x"a6",x"c4"),
  1559 => (x"87",x"d8",x"e0",x"78"),
  1560 => (x"cc",x"48",x"7e",x"70"),
  1561 => (x"c5",x"06",x"a8",x"66"),
  1562 => (x"48",x"a6",x"cc",x"87"),
  1563 => (x"dd",x"ff",x"78",x"6e"),
  1564 => (x"4c",x"70",x"87",x"df"),
  1565 => (x"05",x"ac",x"ec",x"c0"),
  1566 => (x"d0",x"87",x"ee",x"c1"),
  1567 => (x"91",x"cc",x"49",x"66"),
  1568 => (x"81",x"66",x"c4",x"c1"),
  1569 => (x"6a",x"4a",x"a1",x"c4"),
  1570 => (x"4a",x"a1",x"c8",x"4d"),
  1571 => (x"d9",x"c1",x"52",x"6e"),
  1572 => (x"dc",x"ff",x"79",x"d5"),
  1573 => (x"4c",x"70",x"87",x"fb"),
  1574 => (x"87",x"d9",x"02",x"9c"),
  1575 => (x"02",x"ac",x"fb",x"c0"),
  1576 => (x"55",x"74",x"87",x"d3"),
  1577 => (x"87",x"e9",x"dc",x"ff"),
  1578 => (x"02",x"9c",x"4c",x"70"),
  1579 => (x"fb",x"c0",x"87",x"c7"),
  1580 => (x"ed",x"ff",x"05",x"ac"),
  1581 => (x"55",x"e0",x"c0",x"87"),
  1582 => (x"c0",x"55",x"c1",x"c2"),
  1583 => (x"e0",x"c0",x"7d",x"97"),
  1584 => (x"66",x"c4",x"48",x"66"),
  1585 => (x"87",x"db",x"05",x"a8"),
  1586 => (x"d4",x"48",x"66",x"d0"),
  1587 => (x"ca",x"04",x"a8",x"66"),
  1588 => (x"48",x"66",x"d0",x"87"),
  1589 => (x"a6",x"d4",x"80",x"c1"),
  1590 => (x"d4",x"87",x"c8",x"58"),
  1591 => (x"88",x"c1",x"48",x"66"),
  1592 => (x"ff",x"58",x"a6",x"d8"),
  1593 => (x"70",x"87",x"ea",x"db"),
  1594 => (x"ac",x"d0",x"c1",x"4c"),
  1595 => (x"dc",x"87",x"c9",x"05"),
  1596 => (x"80",x"c1",x"48",x"66"),
  1597 => (x"58",x"a6",x"e0",x"c0"),
  1598 => (x"02",x"ac",x"d0",x"c1"),
  1599 => (x"6e",x"87",x"d9",x"fd"),
  1600 => (x"66",x"e0",x"c0",x"48"),
  1601 => (x"ea",x"c9",x"05",x"a8"),
  1602 => (x"a6",x"e4",x"c0",x"87"),
  1603 => (x"74",x"78",x"c0",x"48"),
  1604 => (x"88",x"fb",x"c0",x"48"),
  1605 => (x"70",x"58",x"a6",x"c8"),
  1606 => (x"dc",x"c9",x"02",x"98"),
  1607 => (x"88",x"cb",x"48",x"87"),
  1608 => (x"70",x"58",x"a6",x"c8"),
  1609 => (x"ce",x"c1",x"02",x"98"),
  1610 => (x"88",x"c9",x"48",x"87"),
  1611 => (x"70",x"58",x"a6",x"c8"),
  1612 => (x"fe",x"c3",x"02",x"98"),
  1613 => (x"88",x"c4",x"48",x"87"),
  1614 => (x"70",x"58",x"a6",x"c8"),
  1615 => (x"87",x"cf",x"02",x"98"),
  1616 => (x"c8",x"88",x"c1",x"48"),
  1617 => (x"98",x"70",x"58",x"a6"),
  1618 => (x"87",x"e7",x"c3",x"02"),
  1619 => (x"c8",x"87",x"db",x"c8"),
  1620 => (x"f0",x"c0",x"48",x"a6"),
  1621 => (x"f8",x"d9",x"ff",x"78"),
  1622 => (x"c0",x"4c",x"70",x"87"),
  1623 => (x"c3",x"02",x"ac",x"ec"),
  1624 => (x"5c",x"a6",x"cc",x"87"),
  1625 => (x"02",x"ac",x"ec",x"c0"),
  1626 => (x"d9",x"ff",x"87",x"cd"),
  1627 => (x"4c",x"70",x"87",x"e3"),
  1628 => (x"05",x"ac",x"ec",x"c0"),
  1629 => (x"c0",x"87",x"f3",x"ff"),
  1630 => (x"c0",x"02",x"ac",x"ec"),
  1631 => (x"d9",x"ff",x"87",x"c4"),
  1632 => (x"1e",x"c0",x"87",x"cf"),
  1633 => (x"66",x"d8",x"1e",x"ca"),
  1634 => (x"c1",x"91",x"cc",x"49"),
  1635 => (x"71",x"48",x"66",x"cc"),
  1636 => (x"58",x"a6",x"cc",x"80"),
  1637 => (x"c4",x"48",x"66",x"c8"),
  1638 => (x"58",x"a6",x"d0",x"80"),
  1639 => (x"49",x"bf",x"66",x"cc"),
  1640 => (x"87",x"e9",x"d9",x"ff"),
  1641 => (x"1e",x"de",x"1e",x"c1"),
  1642 => (x"49",x"bf",x"66",x"d4"),
  1643 => (x"87",x"dd",x"d9",x"ff"),
  1644 => (x"49",x"70",x"86",x"d0"),
  1645 => (x"88",x"08",x"c0",x"48"),
  1646 => (x"58",x"a6",x"ec",x"c0"),
  1647 => (x"c0",x"06",x"a8",x"c0"),
  1648 => (x"e8",x"c0",x"87",x"ee"),
  1649 => (x"a8",x"dd",x"48",x"66"),
  1650 => (x"87",x"e4",x"c0",x"03"),
  1651 => (x"49",x"bf",x"66",x"c4"),
  1652 => (x"81",x"66",x"e8",x"c0"),
  1653 => (x"c0",x"51",x"e0",x"c0"),
  1654 => (x"c1",x"49",x"66",x"e8"),
  1655 => (x"bf",x"66",x"c4",x"81"),
  1656 => (x"51",x"c1",x"c2",x"81"),
  1657 => (x"49",x"66",x"e8",x"c0"),
  1658 => (x"66",x"c4",x"81",x"c2"),
  1659 => (x"51",x"c0",x"81",x"bf"),
  1660 => (x"d8",x"c1",x"48",x"6e"),
  1661 => (x"49",x"6e",x"78",x"cf"),
  1662 => (x"66",x"d8",x"81",x"c8"),
  1663 => (x"c9",x"49",x"6e",x"51"),
  1664 => (x"51",x"66",x"dc",x"81"),
  1665 => (x"81",x"ca",x"49",x"6e"),
  1666 => (x"d8",x"51",x"66",x"c8"),
  1667 => (x"80",x"c1",x"48",x"66"),
  1668 => (x"d0",x"58",x"a6",x"dc"),
  1669 => (x"66",x"d4",x"48",x"66"),
  1670 => (x"cb",x"c0",x"04",x"a8"),
  1671 => (x"48",x"66",x"d0",x"87"),
  1672 => (x"a6",x"d4",x"80",x"c1"),
  1673 => (x"87",x"d1",x"c5",x"58"),
  1674 => (x"c1",x"48",x"66",x"d4"),
  1675 => (x"58",x"a6",x"d8",x"88"),
  1676 => (x"ff",x"87",x"c6",x"c5"),
  1677 => (x"c0",x"87",x"c1",x"d9"),
  1678 => (x"ff",x"58",x"a6",x"ec"),
  1679 => (x"c0",x"87",x"f9",x"d8"),
  1680 => (x"c0",x"58",x"a6",x"f0"),
  1681 => (x"c0",x"05",x"a8",x"ec"),
  1682 => (x"48",x"a6",x"87",x"c9"),
  1683 => (x"78",x"66",x"e8",x"c0"),
  1684 => (x"ff",x"87",x"c4",x"c0"),
  1685 => (x"d0",x"87",x"fa",x"d5"),
  1686 => (x"91",x"cc",x"49",x"66"),
  1687 => (x"48",x"66",x"c4",x"c1"),
  1688 => (x"a6",x"c8",x"80",x"71"),
  1689 => (x"4a",x"66",x"c4",x"58"),
  1690 => (x"66",x"c4",x"82",x"c8"),
  1691 => (x"c0",x"81",x"ca",x"49"),
  1692 => (x"c0",x"51",x"66",x"e8"),
  1693 => (x"c1",x"49",x"66",x"ec"),
  1694 => (x"66",x"e8",x"c0",x"81"),
  1695 => (x"71",x"48",x"c1",x"89"),
  1696 => (x"c1",x"49",x"70",x"30"),
  1697 => (x"7a",x"97",x"71",x"89"),
  1698 => (x"bf",x"c8",x"f7",x"c2"),
  1699 => (x"66",x"e8",x"c0",x"49"),
  1700 => (x"4a",x"6a",x"97",x"29"),
  1701 => (x"c0",x"98",x"71",x"48"),
  1702 => (x"c4",x"58",x"a6",x"f4"),
  1703 => (x"80",x"c4",x"48",x"66"),
  1704 => (x"c8",x"58",x"a6",x"cc"),
  1705 => (x"c0",x"4d",x"bf",x"66"),
  1706 => (x"6e",x"48",x"66",x"e0"),
  1707 => (x"c5",x"c0",x"02",x"a8"),
  1708 => (x"c0",x"7e",x"c0",x"87"),
  1709 => (x"7e",x"c1",x"87",x"c2"),
  1710 => (x"e0",x"c0",x"1e",x"6e"),
  1711 => (x"ff",x"49",x"75",x"1e"),
  1712 => (x"c8",x"87",x"ca",x"d5"),
  1713 => (x"c0",x"4c",x"70",x"86"),
  1714 => (x"c1",x"06",x"ac",x"b7"),
  1715 => (x"85",x"74",x"87",x"d4"),
  1716 => (x"49",x"bf",x"66",x"c8"),
  1717 => (x"75",x"81",x"e0",x"c0"),
  1718 => (x"f0",x"c1",x"4b",x"89"),
  1719 => (x"fe",x"71",x"4a",x"e8"),
  1720 => (x"c2",x"87",x"c1",x"d9"),
  1721 => (x"c0",x"7e",x"75",x"85"),
  1722 => (x"c1",x"48",x"66",x"e4"),
  1723 => (x"a6",x"e8",x"c0",x"80"),
  1724 => (x"66",x"f0",x"c0",x"58"),
  1725 => (x"70",x"81",x"c1",x"49"),
  1726 => (x"c5",x"c0",x"02",x"a9"),
  1727 => (x"c0",x"4d",x"c0",x"87"),
  1728 => (x"4d",x"c1",x"87",x"c2"),
  1729 => (x"66",x"cc",x"1e",x"75"),
  1730 => (x"e0",x"c0",x"49",x"bf"),
  1731 => (x"89",x"66",x"c4",x"81"),
  1732 => (x"66",x"c8",x"1e",x"71"),
  1733 => (x"f4",x"d3",x"ff",x"49"),
  1734 => (x"c0",x"86",x"c8",x"87"),
  1735 => (x"ff",x"01",x"a8",x"b7"),
  1736 => (x"e4",x"c0",x"87",x"c5"),
  1737 => (x"d3",x"c0",x"02",x"66"),
  1738 => (x"49",x"66",x"c4",x"87"),
  1739 => (x"e4",x"c0",x"81",x"c9"),
  1740 => (x"66",x"c4",x"51",x"66"),
  1741 => (x"e3",x"da",x"c1",x"48"),
  1742 => (x"87",x"ce",x"c0",x"78"),
  1743 => (x"c9",x"49",x"66",x"c4"),
  1744 => (x"c4",x"51",x"c2",x"81"),
  1745 => (x"dc",x"c1",x"48",x"66"),
  1746 => (x"66",x"d0",x"78",x"e1"),
  1747 => (x"a8",x"66",x"d4",x"48"),
  1748 => (x"87",x"cb",x"c0",x"04"),
  1749 => (x"c1",x"48",x"66",x"d0"),
  1750 => (x"58",x"a6",x"d4",x"80"),
  1751 => (x"d4",x"87",x"da",x"c0"),
  1752 => (x"88",x"c1",x"48",x"66"),
  1753 => (x"c0",x"58",x"a6",x"d8"),
  1754 => (x"d2",x"ff",x"87",x"cf"),
  1755 => (x"4c",x"70",x"87",x"cb"),
  1756 => (x"ff",x"87",x"c6",x"c0"),
  1757 => (x"70",x"87",x"c2",x"d2"),
  1758 => (x"48",x"66",x"dc",x"4c"),
  1759 => (x"e0",x"c0",x"80",x"c1"),
  1760 => (x"9c",x"74",x"58",x"a6"),
  1761 => (x"87",x"cb",x"c0",x"02"),
  1762 => (x"c1",x"48",x"66",x"d0"),
  1763 => (x"04",x"a8",x"66",x"cc"),
  1764 => (x"d0",x"87",x"f2",x"f2"),
  1765 => (x"a8",x"c7",x"48",x"66"),
  1766 => (x"87",x"e1",x"c0",x"03"),
  1767 => (x"c2",x"4c",x"66",x"d0"),
  1768 => (x"c0",x"48",x"e0",x"f8"),
  1769 => (x"cc",x"49",x"74",x"78"),
  1770 => (x"66",x"c4",x"c1",x"91"),
  1771 => (x"4a",x"a1",x"c4",x"81"),
  1772 => (x"52",x"c0",x"4a",x"6a"),
  1773 => (x"c7",x"84",x"c1",x"79"),
  1774 => (x"e2",x"ff",x"04",x"ac"),
  1775 => (x"66",x"e0",x"c0",x"87"),
  1776 => (x"87",x"e2",x"c0",x"02"),
  1777 => (x"49",x"66",x"c4",x"c1"),
  1778 => (x"c1",x"81",x"d4",x"c1"),
  1779 => (x"c1",x"4a",x"66",x"c4"),
  1780 => (x"52",x"c0",x"82",x"dc"),
  1781 => (x"79",x"d5",x"d9",x"c1"),
  1782 => (x"49",x"66",x"c4",x"c1"),
  1783 => (x"c1",x"81",x"d8",x"c1"),
  1784 => (x"c0",x"79",x"ec",x"f0"),
  1785 => (x"c4",x"c1",x"87",x"d6"),
  1786 => (x"d4",x"c1",x"49",x"66"),
  1787 => (x"66",x"c4",x"c1",x"81"),
  1788 => (x"82",x"d8",x"c1",x"4a"),
  1789 => (x"7a",x"f4",x"f0",x"c1"),
  1790 => (x"79",x"cc",x"d9",x"c1"),
  1791 => (x"49",x"66",x"c4",x"c1"),
  1792 => (x"c1",x"81",x"e0",x"c1"),
  1793 => (x"ff",x"79",x"f3",x"dc"),
  1794 => (x"cc",x"87",x"e5",x"cf"),
  1795 => (x"cc",x"ff",x"48",x"66"),
  1796 => (x"26",x"4d",x"26",x"8e"),
  1797 => (x"26",x"4b",x"26",x"4c"),
  1798 => (x"00",x"00",x"00",x"4f"),
  1799 => (x"64",x"61",x"6f",x"4c"),
  1800 => (x"20",x"2e",x"2a",x"20"),
  1801 => (x"00",x"00",x"00",x"00"),
  1802 => (x"00",x"00",x"20",x"3a"),
  1803 => (x"61",x"42",x"20",x"80"),
  1804 => (x"00",x"00",x"6b",x"63"),
  1805 => (x"78",x"45",x"20",x"80"),
  1806 => (x"1e",x"00",x"74",x"69"),
  1807 => (x"f8",x"c2",x"1e",x"c7"),
  1808 => (x"c1",x"1e",x"bf",x"dc"),
  1809 => (x"c2",x"1e",x"cc",x"f4"),
  1810 => (x"bf",x"97",x"cc",x"f7"),
  1811 => (x"87",x"f5",x"ec",x"49"),
  1812 => (x"49",x"cc",x"f4",x"c1"),
  1813 => (x"87",x"e6",x"e2",x"c0"),
  1814 => (x"4f",x"26",x"8e",x"f4"),
  1815 => (x"c8",x"1e",x"73",x"1e"),
  1816 => (x"f5",x"c1",x"87",x"c3"),
  1817 => (x"f3",x"c1",x"48",x"e4"),
  1818 => (x"e8",x"fe",x"78",x"ec"),
  1819 => (x"e2",x"c0",x"49",x"a0"),
  1820 => (x"49",x"c7",x"87",x"cc"),
  1821 => (x"87",x"f8",x"e0",x"c0"),
  1822 => (x"e2",x"c0",x"49",x"c1"),
  1823 => (x"d4",x"ff",x"87",x"d3"),
  1824 => (x"78",x"ff",x"c3",x"48"),
  1825 => (x"48",x"e8",x"f8",x"c2"),
  1826 => (x"dd",x"fe",x"50",x"c0"),
  1827 => (x"98",x"70",x"87",x"e2"),
  1828 => (x"fe",x"87",x"cd",x"02"),
  1829 => (x"70",x"87",x"de",x"e7"),
  1830 => (x"87",x"c4",x"02",x"98"),
  1831 => (x"87",x"c2",x"4a",x"c1"),
  1832 => (x"9a",x"72",x"4a",x"c0"),
  1833 => (x"c1",x"87",x"c8",x"02"),
  1834 => (x"fe",x"49",x"f8",x"f3"),
  1835 => (x"c2",x"87",x"f8",x"cf"),
  1836 => (x"c0",x"48",x"dc",x"f8"),
  1837 => (x"cc",x"f7",x"c2",x"78"),
  1838 => (x"49",x"50",x"c0",x"48"),
  1839 => (x"c0",x"87",x"fc",x"fd"),
  1840 => (x"70",x"87",x"ea",x"f5"),
  1841 => (x"cb",x"02",x"9b",x"4b"),
  1842 => (x"e8",x"f5",x"c1",x"87"),
  1843 => (x"df",x"49",x"c7",x"5b"),
  1844 => (x"87",x"c6",x"87",x"de"),
  1845 => (x"e0",x"c0",x"49",x"c0"),
  1846 => (x"c2",x"c3",x"87",x"f7"),
  1847 => (x"d8",x"e2",x"c0",x"87"),
  1848 => (x"ec",x"ef",x"c0",x"87"),
  1849 => (x"87",x"f5",x"ff",x"87"),
  1850 => (x"4f",x"26",x"4b",x"26"),
  1851 => (x"74",x"6f",x"6f",x"42"),
  1852 => (x"2e",x"67",x"6e",x"69"),
  1853 => (x"00",x"00",x"2e",x"2e"),
  1854 => (x"4f",x"20",x"44",x"53"),
  1855 => (x"00",x"00",x"00",x"4b"),
  1856 => (x"00",x"00",x"00",x"00"),
  1857 => (x"00",x"00",x"00",x"00"),
  1858 => (x"00",x"00",x"00",x"01"),
  1859 => (x"00",x"00",x"13",x"3b"),
  1860 => (x"00",x"00",x"2e",x"34"),
  1861 => (x"00",x"00",x"00",x"00"),
  1862 => (x"00",x"00",x"13",x"3b"),
  1863 => (x"00",x"00",x"2e",x"52"),
  1864 => (x"00",x"00",x"00",x"00"),
  1865 => (x"00",x"00",x"13",x"3b"),
  1866 => (x"00",x"00",x"2e",x"70"),
  1867 => (x"00",x"00",x"00",x"00"),
  1868 => (x"00",x"00",x"13",x"3b"),
  1869 => (x"00",x"00",x"2e",x"8e"),
  1870 => (x"00",x"00",x"00",x"00"),
  1871 => (x"00",x"00",x"13",x"3b"),
  1872 => (x"00",x"00",x"2e",x"ac"),
  1873 => (x"00",x"00",x"00",x"00"),
  1874 => (x"00",x"00",x"13",x"3b"),
  1875 => (x"00",x"00",x"2e",x"ca"),
  1876 => (x"00",x"00",x"00",x"00"),
  1877 => (x"00",x"00",x"13",x"3b"),
  1878 => (x"00",x"00",x"2e",x"e8"),
  1879 => (x"00",x"00",x"00",x"00"),
  1880 => (x"00",x"00",x"16",x"55"),
  1881 => (x"00",x"00",x"00",x"00"),
  1882 => (x"00",x"00",x"00",x"00"),
  1883 => (x"00",x"00",x"13",x"ef"),
  1884 => (x"00",x"00",x"00",x"00"),
  1885 => (x"00",x"00",x"00",x"00"),
  1886 => (x"db",x"86",x"fc",x"1e"),
  1887 => (x"fc",x"7e",x"70",x"87"),
  1888 => (x"1e",x"4f",x"26",x"8e"),
  1889 => (x"c0",x"48",x"f0",x"fe"),
  1890 => (x"79",x"09",x"cd",x"78"),
  1891 => (x"1e",x"4f",x"26",x"09"),
  1892 => (x"49",x"f8",x"f5",x"c1"),
  1893 => (x"4f",x"26",x"87",x"ed"),
  1894 => (x"bf",x"f0",x"fe",x"1e"),
  1895 => (x"1e",x"4f",x"26",x"48"),
  1896 => (x"c1",x"48",x"f0",x"fe"),
  1897 => (x"1e",x"4f",x"26",x"78"),
  1898 => (x"c0",x"48",x"f0",x"fe"),
  1899 => (x"1e",x"4f",x"26",x"78"),
  1900 => (x"52",x"c0",x"4a",x"71"),
  1901 => (x"0e",x"4f",x"26",x"51"),
  1902 => (x"5d",x"5c",x"5b",x"5e"),
  1903 => (x"71",x"86",x"f4",x"0e"),
  1904 => (x"7e",x"6d",x"97",x"4d"),
  1905 => (x"97",x"4c",x"a5",x"c1"),
  1906 => (x"a6",x"c8",x"48",x"6c"),
  1907 => (x"c4",x"48",x"6e",x"58"),
  1908 => (x"c5",x"05",x"a8",x"66"),
  1909 => (x"c0",x"48",x"ff",x"87"),
  1910 => (x"ca",x"ff",x"87",x"e6"),
  1911 => (x"49",x"a5",x"c2",x"87"),
  1912 => (x"71",x"4b",x"6c",x"97"),
  1913 => (x"6b",x"97",x"4b",x"a3"),
  1914 => (x"7e",x"6c",x"97",x"4b"),
  1915 => (x"80",x"c1",x"48",x"6e"),
  1916 => (x"c7",x"58",x"a6",x"c8"),
  1917 => (x"58",x"a6",x"cc",x"98"),
  1918 => (x"fe",x"7c",x"97",x"70"),
  1919 => (x"48",x"73",x"87",x"e1"),
  1920 => (x"4d",x"26",x"8e",x"f4"),
  1921 => (x"4b",x"26",x"4c",x"26"),
  1922 => (x"5e",x"0e",x"4f",x"26"),
  1923 => (x"f4",x"0e",x"5c",x"5b"),
  1924 => (x"d8",x"4c",x"71",x"86"),
  1925 => (x"ff",x"c3",x"4a",x"66"),
  1926 => (x"4b",x"a4",x"c2",x"9a"),
  1927 => (x"73",x"49",x"6c",x"97"),
  1928 => (x"51",x"72",x"49",x"a1"),
  1929 => (x"6e",x"7e",x"6c",x"97"),
  1930 => (x"c8",x"80",x"c1",x"48"),
  1931 => (x"98",x"c7",x"58",x"a6"),
  1932 => (x"70",x"58",x"a6",x"cc"),
  1933 => (x"26",x"8e",x"f4",x"54"),
  1934 => (x"26",x"4b",x"26",x"4c"),
  1935 => (x"86",x"fc",x"1e",x"4f"),
  1936 => (x"e0",x"87",x"e4",x"fd"),
  1937 => (x"c0",x"49",x"4a",x"bf"),
  1938 => (x"02",x"99",x"c0",x"e0"),
  1939 => (x"1e",x"72",x"87",x"cb"),
  1940 => (x"49",x"c8",x"fc",x"c2"),
  1941 => (x"c4",x"87",x"f3",x"fe"),
  1942 => (x"87",x"fc",x"fc",x"86"),
  1943 => (x"fe",x"fc",x"7e",x"70"),
  1944 => (x"26",x"8e",x"fc",x"87"),
  1945 => (x"fc",x"c2",x"1e",x"4f"),
  1946 => (x"c2",x"fd",x"49",x"c8"),
  1947 => (x"fd",x"f8",x"c1",x"87"),
  1948 => (x"87",x"cf",x"fc",x"49"),
  1949 => (x"26",x"87",x"ed",x"c3"),
  1950 => (x"5b",x"5e",x"0e",x"4f"),
  1951 => (x"fc",x"0e",x"5d",x"5c"),
  1952 => (x"ff",x"7e",x"71",x"86"),
  1953 => (x"fc",x"c2",x"4d",x"d4"),
  1954 => (x"ea",x"fc",x"49",x"c8"),
  1955 => (x"c0",x"4b",x"70",x"87"),
  1956 => (x"c2",x"04",x"ab",x"b7"),
  1957 => (x"f0",x"c3",x"87",x"f8"),
  1958 => (x"87",x"c9",x"05",x"ab"),
  1959 => (x"48",x"dc",x"fd",x"c1"),
  1960 => (x"d9",x"c2",x"78",x"c1"),
  1961 => (x"ab",x"e0",x"c3",x"87"),
  1962 => (x"c1",x"87",x"c9",x"05"),
  1963 => (x"c1",x"48",x"e0",x"fd"),
  1964 => (x"87",x"ca",x"c2",x"78"),
  1965 => (x"bf",x"e0",x"fd",x"c1"),
  1966 => (x"c2",x"87",x"c6",x"02"),
  1967 => (x"c2",x"4c",x"a3",x"c0"),
  1968 => (x"c1",x"4c",x"73",x"87"),
  1969 => (x"02",x"bf",x"dc",x"fd"),
  1970 => (x"74",x"87",x"e0",x"c0"),
  1971 => (x"29",x"b7",x"c4",x"49"),
  1972 => (x"f8",x"fe",x"c1",x"91"),
  1973 => (x"cf",x"4a",x"74",x"81"),
  1974 => (x"c1",x"92",x"c2",x"9a"),
  1975 => (x"70",x"30",x"72",x"48"),
  1976 => (x"72",x"ba",x"ff",x"4a"),
  1977 => (x"70",x"98",x"69",x"48"),
  1978 => (x"74",x"87",x"db",x"79"),
  1979 => (x"29",x"b7",x"c4",x"49"),
  1980 => (x"f8",x"fe",x"c1",x"91"),
  1981 => (x"cf",x"4a",x"74",x"81"),
  1982 => (x"c3",x"92",x"c2",x"9a"),
  1983 => (x"70",x"30",x"72",x"48"),
  1984 => (x"b0",x"69",x"48",x"4a"),
  1985 => (x"05",x"6e",x"79",x"70"),
  1986 => (x"ff",x"87",x"e7",x"c0"),
  1987 => (x"e1",x"c8",x"48",x"d0"),
  1988 => (x"c1",x"7d",x"c5",x"78"),
  1989 => (x"02",x"bf",x"e0",x"fd"),
  1990 => (x"e0",x"c3",x"87",x"c3"),
  1991 => (x"dc",x"fd",x"c1",x"7d"),
  1992 => (x"87",x"c3",x"02",x"bf"),
  1993 => (x"73",x"7d",x"f0",x"c3"),
  1994 => (x"48",x"d0",x"ff",x"7d"),
  1995 => (x"c0",x"78",x"e1",x"c8"),
  1996 => (x"fd",x"c1",x"78",x"e0"),
  1997 => (x"78",x"c0",x"48",x"e0"),
  1998 => (x"48",x"dc",x"fd",x"c1"),
  1999 => (x"fc",x"c2",x"78",x"c0"),
  2000 => (x"f2",x"f9",x"49",x"c8"),
  2001 => (x"c0",x"4b",x"70",x"87"),
  2002 => (x"fd",x"03",x"ab",x"b7"),
  2003 => (x"48",x"c0",x"87",x"c8"),
  2004 => (x"4d",x"26",x"8e",x"fc"),
  2005 => (x"4b",x"26",x"4c",x"26"),
  2006 => (x"00",x"00",x"4f",x"26"),
  2007 => (x"00",x"00",x"00",x"00"),
  2008 => (x"00",x"00",x"00",x"00"),
  2009 => (x"72",x"4a",x"c0",x"1e"),
  2010 => (x"c1",x"91",x"c4",x"49"),
  2011 => (x"c0",x"81",x"f8",x"fe"),
  2012 => (x"d0",x"82",x"c1",x"79"),
  2013 => (x"ee",x"04",x"aa",x"b7"),
  2014 => (x"0e",x"4f",x"26",x"87"),
  2015 => (x"5d",x"5c",x"5b",x"5e"),
  2016 => (x"f8",x"4d",x"71",x"0e"),
  2017 => (x"4a",x"75",x"87",x"e1"),
  2018 => (x"92",x"2a",x"b7",x"c4"),
  2019 => (x"82",x"f8",x"fe",x"c1"),
  2020 => (x"9c",x"cf",x"4c",x"75"),
  2021 => (x"49",x"6a",x"94",x"c2"),
  2022 => (x"c3",x"2b",x"74",x"4b"),
  2023 => (x"74",x"48",x"c2",x"9b"),
  2024 => (x"ff",x"4c",x"70",x"30"),
  2025 => (x"71",x"48",x"74",x"bc"),
  2026 => (x"f7",x"7a",x"70",x"98"),
  2027 => (x"48",x"73",x"87",x"f1"),
  2028 => (x"4c",x"26",x"4d",x"26"),
  2029 => (x"4f",x"26",x"4b",x"26"),
  2030 => (x"00",x"00",x"00",x"00"),
  2031 => (x"00",x"00",x"00",x"00"),
  2032 => (x"00",x"00",x"00",x"00"),
  2033 => (x"00",x"00",x"00",x"00"),
  2034 => (x"00",x"00",x"00",x"00"),
  2035 => (x"00",x"00",x"00",x"00"),
  2036 => (x"00",x"00",x"00",x"00"),
  2037 => (x"00",x"00",x"00",x"00"),
  2038 => (x"00",x"00",x"00",x"00"),
  2039 => (x"00",x"00",x"00",x"00"),
  2040 => (x"00",x"00",x"00",x"00"),
  2041 => (x"00",x"00",x"00",x"00"),
  2042 => (x"00",x"00",x"00",x"00"),
  2043 => (x"00",x"00",x"00",x"00"),
  2044 => (x"00",x"00",x"00",x"00"),
  2045 => (x"00",x"00",x"00",x"00"),
  2046 => (x"48",x"d0",x"ff",x"1e"),
  2047 => (x"71",x"78",x"e1",x"c8"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

